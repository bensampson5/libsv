module decoder_8b10b (
    input  logic [9:0] i_10b,
    input  logic       i_disp,
    output logic [7:0] o_8b,
    output logic       o_disp,
    output logic       o_ctrl,
    output logic       o_code_err,
    output logic       o_disp_err
);

  // Placeholder implementation for testbench development (will fail)
  assign o_8b       = '0;
  assign o_disp     = '0;
  assign o_ctrl     = '0;
  assign o_code_err = '0;
  assign o_disp_err = '0;

endmodule
