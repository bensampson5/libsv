module encoder_8b10b (
    input  logic [7:0] i_8b,
    input  logic       i_rd,
    input  logic       i_ctrl,
    output logic [9:0] o_10b,
    output logic       o_rd
);

  // Create lookup table input and output vectors
  logic [ 9:0] i_lut;
  logic [10:0] o_lut;
  assign i_lut = {i_ctrl, i_rd, i_8b};
  assign o_rd  = o_lut[10];
  assign o_10b = o_lut[9:0];

  // Mapping is XRHGFEDCBA: rjhgfiedcba, where X selects a control symbol if
  // '1', R is the input running disparity (0 = -1, 1 = +1), and r is the
  // output running disparity (0 = -1, 1 = +1)
  always_comb begin
    case (i_lut)
      //  XRHGFEDCBA:             rjhgfiedbca
      10'b0000000000: o_lut = 11'b00010111001;  // D.00.0, RDin = -1, RDout = -1
      10'b0000000001: o_lut = 11'b00010101110;  // D.01.0, RDin = -1, RDout = -1
      10'b0000000010: o_lut = 11'b00010101101;  // D.02.0, RDin = -1, RDout = -1
      10'b0000000011: o_lut = 11'b11101100011;  // D.03.0, RDin = -1, RDout = +1
      10'b0000000100: o_lut = 11'b00010101011;  // D.04.0, RDin = -1, RDout = -1
      10'b0000000101: o_lut = 11'b11101100101;  // D.05.0, RDin = -1, RDout = +1
      10'b0000000110: o_lut = 11'b11101100110;  // D.06.0, RDin = -1, RDout = +1
      10'b0000000111: o_lut = 11'b11101000111;  // D.07.0, RDin = -1, RDout = +1
      10'b0000001000: o_lut = 11'b00010100111;  // D.08.0, RDin = -1, RDout = -1
      10'b0000001001: o_lut = 11'b11101101001;  // D.09.0, RDin = -1, RDout = +1
      10'b0000001010: o_lut = 11'b11101101010;  // D.10.0, RDin = -1, RDout = +1
      10'b0000001011: o_lut = 11'b11101001011;  // D.11.0, RDin = -1, RDout = +1
      10'b0000001100: o_lut = 11'b11101101100;  // D.12.0, RDin = -1, RDout = +1
      10'b0000001101: o_lut = 11'b11101001101;  // D.13.0, RDin = -1, RDout = +1
      10'b0000001110: o_lut = 11'b11101001110;  // D.14.0, RDin = -1, RDout = +1
      10'b0000001111: o_lut = 11'b00010111010;  // D.15.0, RDin = -1, RDout = -1
      10'b0000010000: o_lut = 11'b00010110110;  // D.16.0, RDin = -1, RDout = -1
      10'b0000010001: o_lut = 11'b11101110001;  // D.17.0, RDin = -1, RDout = +1
      10'b0000010010: o_lut = 11'b11101110010;  // D.18.0, RDin = -1, RDout = +1
      10'b0000010011: o_lut = 11'b11101010011;  // D.19.0, RDin = -1, RDout = +1
      10'b0000010100: o_lut = 11'b11101110100;  // D.20.0, RDin = -1, RDout = +1
      10'b0000010101: o_lut = 11'b11101010101;  // D.21.0, RDin = -1, RDout = +1
      10'b0000010110: o_lut = 11'b11101010110;  // D.22.0, RDin = -1, RDout = +1
      10'b0000010111: o_lut = 11'b00010010111;  // D.23.0, RDin = -1, RDout = -1
      10'b0000011000: o_lut = 11'b00010110011;  // D.24.0, RDin = -1, RDout = -1
      10'b0000011001: o_lut = 11'b11101011001;  // D.25.0, RDin = -1, RDout = +1
      10'b0000011010: o_lut = 11'b11101011010;  // D.26.0, RDin = -1, RDout = +1
      10'b0000011011: o_lut = 11'b00010011011;  // D.27.0, RDin = -1, RDout = -1
      10'b0000011100: o_lut = 11'b11101001110;  // D.28.0, RDin = -1, RDout = +1
      10'b0000011101: o_lut = 11'b00010011101;  // D.29.0, RDin = -1, RDout = -1
      10'b0000011110: o_lut = 11'b00010011110;  // D.30.0, RDin = -1, RDout = -1
      10'b0000011111: o_lut = 11'b00010110101;  // D.31.0, RDin = -1, RDout = -1
      10'b0000100000: o_lut = 11'b11001111001;  // D.00.1, RDin = -1, RDout = +1
      10'b0000100001: o_lut = 11'b11001101110;  // D.01.1, RDin = -1, RDout = +1
      10'b0000100010: o_lut = 11'b11001101101;  // D.02.1, RDin = -1, RDout = +1
      10'b0000100011: o_lut = 11'b01001100011;  // D.03.1, RDin = -1, RDout = -1
      10'b0000100100: o_lut = 11'b11001101011;  // D.04.1, RDin = -1, RDout = +1
      10'b0000100101: o_lut = 11'b01001100101;  // D.05.1, RDin = -1, RDout = -1
      10'b0000100110: o_lut = 11'b01001100110;  // D.06.1, RDin = -1, RDout = -1
      10'b0000100111: o_lut = 11'b01001000111;  // D.07.1, RDin = -1, RDout = -1
      10'b0000101000: o_lut = 11'b11001100111;  // D.08.1, RDin = -1, RDout = +1
      10'b0000101001: o_lut = 11'b01001101001;  // D.09.1, RDin = -1, RDout = -1
      10'b0000101010: o_lut = 11'b01001101010;  // D.10.1, RDin = -1, RDout = -1
      10'b0000101011: o_lut = 11'b01001001011;  // D.11.1, RDin = -1, RDout = -1
      10'b0000101100: o_lut = 11'b01001101100;  // D.12.1, RDin = -1, RDout = -1
      10'b0000101101: o_lut = 11'b01001001101;  // D.13.1, RDin = -1, RDout = -1
      10'b0000101110: o_lut = 11'b01001001110;  // D.14.1, RDin = -1, RDout = -1
      10'b0000101111: o_lut = 11'b11001111010;  // D.15.1, RDin = -1, RDout = +1
      10'b0000110000: o_lut = 11'b11001110110;  // D.16.1, RDin = -1, RDout = +1
      10'b0000110001: o_lut = 11'b01001110001;  // D.17.1, RDin = -1, RDout = -1
      10'b0000110010: o_lut = 11'b01001110010;  // D.18.1, RDin = -1, RDout = -1
      10'b0000110011: o_lut = 11'b01001010011;  // D.19.1, RDin = -1, RDout = -1
      10'b0000110100: o_lut = 11'b01001110100;  // D.20.1, RDin = -1, RDout = -1
      10'b0000110101: o_lut = 11'b01001010101;  // D.21.1, RDin = -1, RDout = -1
      10'b0000110110: o_lut = 11'b01001010110;  // D.22.1, RDin = -1, RDout = -1
      10'b0000110111: o_lut = 11'b11001010111;  // D.23.1, RDin = -1, RDout = +1
      10'b0000111000: o_lut = 11'b11001110011;  // D.24.1, RDin = -1, RDout = +1
      10'b0000111001: o_lut = 11'b01001011001;  // D.25.1, RDin = -1, RDout = -1
      10'b0000111010: o_lut = 11'b01001011010;  // D.26.1, RDin = -1, RDout = -1
      10'b0000111011: o_lut = 11'b11001011011;  // D.27.1, RDin = -1, RDout = +1
      10'b0000111100: o_lut = 11'b01001001110;  // D.28.1, RDin = -1, RDout = -1
      10'b0000111101: o_lut = 11'b11001011101;  // D.29.1, RDin = -1, RDout = +1
      10'b0000111110: o_lut = 11'b11001011110;  // D.30.1, RDin = -1, RDout = +1
      10'b0000111111: o_lut = 11'b11001110101;  // D.31.1, RDin = -1, RDout = +1
      10'b0001000000: o_lut = 11'b11010111001;  // D.00.2, RDin = -1, RDout = +1
      10'b0001000001: o_lut = 11'b11010101110;  // D.01.2, RDin = -1, RDout = +1
      10'b0001000010: o_lut = 11'b11010101101;  // D.02.2, RDin = -1, RDout = +1
      10'b0001000011: o_lut = 11'b01010100011;  // D.03.2, RDin = -1, RDout = -1
      10'b0001000100: o_lut = 11'b11010101011;  // D.04.2, RDin = -1, RDout = +1
      10'b0001000101: o_lut = 11'b01010100101;  // D.05.2, RDin = -1, RDout = -1
      10'b0001000110: o_lut = 11'b01010100110;  // D.06.2, RDin = -1, RDout = -1
      10'b0001000111: o_lut = 11'b01010000111;  // D.07.2, RDin = -1, RDout = -1
      10'b0001001000: o_lut = 11'b11010100111;  // D.08.2, RDin = -1, RDout = +1
      10'b0001001001: o_lut = 11'b01010101001;  // D.09.2, RDin = -1, RDout = -1
      10'b0001001010: o_lut = 11'b01010101010;  // D.10.2, RDin = -1, RDout = -1
      10'b0001001011: o_lut = 11'b01010001011;  // D.11.2, RDin = -1, RDout = -1
      10'b0001001100: o_lut = 11'b01010101100;  // D.12.2, RDin = -1, RDout = -1
      10'b0001001101: o_lut = 11'b01010001101;  // D.13.2, RDin = -1, RDout = -1
      10'b0001001110: o_lut = 11'b01010001110;  // D.14.2, RDin = -1, RDout = -1
      10'b0001001111: o_lut = 11'b11010111010;  // D.15.2, RDin = -1, RDout = +1
      10'b0001010000: o_lut = 11'b11010110110;  // D.16.2, RDin = -1, RDout = +1
      10'b0001010001: o_lut = 11'b01010110001;  // D.17.2, RDin = -1, RDout = -1
      10'b0001010010: o_lut = 11'b01010110010;  // D.18.2, RDin = -1, RDout = -1
      10'b0001010011: o_lut = 11'b01010010011;  // D.19.2, RDin = -1, RDout = -1
      10'b0001010100: o_lut = 11'b01010110100;  // D.20.2, RDin = -1, RDout = -1
      10'b0001010101: o_lut = 11'b01010010101;  // D.21.2, RDin = -1, RDout = -1
      10'b0001010110: o_lut = 11'b01010010110;  // D.22.2, RDin = -1, RDout = -1
      10'b0001010111: o_lut = 11'b11010010111;  // D.23.2, RDin = -1, RDout = +1
      10'b0001011000: o_lut = 11'b11010110011;  // D.24.2, RDin = -1, RDout = +1
      10'b0001011001: o_lut = 11'b01010011001;  // D.25.2, RDin = -1, RDout = -1
      10'b0001011010: o_lut = 11'b01010011010;  // D.26.2, RDin = -1, RDout = -1
      10'b0001011011: o_lut = 11'b11010011011;  // D.27.2, RDin = -1, RDout = +1
      10'b0001011100: o_lut = 11'b01010001110;  // D.28.2, RDin = -1, RDout = -1
      10'b0001011101: o_lut = 11'b11010011101;  // D.29.2, RDin = -1, RDout = +1
      10'b0001011110: o_lut = 11'b11010011110;  // D.30.2, RDin = -1, RDout = +1
      10'b0001011111: o_lut = 11'b11010110101;  // D.31.2, RDin = -1, RDout = +1
      10'b0001100000: o_lut = 11'b11100111001;  // D.00.3, RDin = -1, RDout = +1
      10'b0001100001: o_lut = 11'b11100101110;  // D.01.3, RDin = -1, RDout = +1
      10'b0001100010: o_lut = 11'b11100101101;  // D.02.3, RDin = -1, RDout = +1
      10'b0001100011: o_lut = 11'b00011100011;  // D.03.3, RDin = -1, RDout = -1
      10'b0001100100: o_lut = 11'b11100101011;  // D.04.3, RDin = -1, RDout = +1
      10'b0001100101: o_lut = 11'b00011100101;  // D.05.3, RDin = -1, RDout = -1
      10'b0001100110: o_lut = 11'b00011100110;  // D.06.3, RDin = -1, RDout = -1
      10'b0001100111: o_lut = 11'b00011000111;  // D.07.3, RDin = -1, RDout = -1
      10'b0001101000: o_lut = 11'b11100100111;  // D.08.3, RDin = -1, RDout = +1
      10'b0001101001: o_lut = 11'b00011101001;  // D.09.3, RDin = -1, RDout = -1
      10'b0001101010: o_lut = 11'b00011101010;  // D.10.3, RDin = -1, RDout = -1
      10'b0001101011: o_lut = 11'b00011001011;  // D.11.3, RDin = -1, RDout = -1
      10'b0001101100: o_lut = 11'b00011101100;  // D.12.3, RDin = -1, RDout = -1
      10'b0001101101: o_lut = 11'b00011001101;  // D.13.3, RDin = -1, RDout = -1
      10'b0001101110: o_lut = 11'b00011001110;  // D.14.3, RDin = -1, RDout = -1
      10'b0001101111: o_lut = 11'b11100111010;  // D.15.3, RDin = -1, RDout = +1
      10'b0001110000: o_lut = 11'b11100110110;  // D.16.3, RDin = -1, RDout = +1
      10'b0001110001: o_lut = 11'b00011110001;  // D.17.3, RDin = -1, RDout = -1
      10'b0001110010: o_lut = 11'b00011110010;  // D.18.3, RDin = -1, RDout = -1
      10'b0001110011: o_lut = 11'b00011010011;  // D.19.3, RDin = -1, RDout = -1
      10'b0001110100: o_lut = 11'b00011110100;  // D.20.3, RDin = -1, RDout = -1
      10'b0001110101: o_lut = 11'b00011010101;  // D.21.3, RDin = -1, RDout = -1
      10'b0001110110: o_lut = 11'b00011010110;  // D.22.3, RDin = -1, RDout = -1
      10'b0001110111: o_lut = 11'b11100010111;  // D.23.3, RDin = -1, RDout = +1
      10'b0001111000: o_lut = 11'b11100110011;  // D.24.3, RDin = -1, RDout = +1
      10'b0001111001: o_lut = 11'b00011011001;  // D.25.3, RDin = -1, RDout = -1
      10'b0001111010: o_lut = 11'b00011011010;  // D.26.3, RDin = -1, RDout = -1
      10'b0001111011: o_lut = 11'b11100011011;  // D.27.3, RDin = -1, RDout = +1
      10'b0001111100: o_lut = 11'b00011001110;  // D.28.3, RDin = -1, RDout = -1
      10'b0001111101: o_lut = 11'b11100011101;  // D.29.3, RDin = -1, RDout = +1
      10'b0001111110: o_lut = 11'b11100011110;  // D.30.3, RDin = -1, RDout = +1
      10'b0001111111: o_lut = 11'b11100110101;  // D.31.3, RDin = -1, RDout = +1
      10'b0010000000: o_lut = 11'b00100111001;  // D.00.4, RDin = -1, RDout = -1
      10'b0010000001: o_lut = 11'b00100101110;  // D.01.4, RDin = -1, RDout = -1
      10'b0010000010: o_lut = 11'b00100101101;  // D.02.4, RDin = -1, RDout = -1
      10'b0010000011: o_lut = 11'b11011100011;  // D.03.4, RDin = -1, RDout = +1
      10'b0010000100: o_lut = 11'b00100101011;  // D.04.4, RDin = -1, RDout = -1
      10'b0010000101: o_lut = 11'b11011100101;  // D.05.4, RDin = -1, RDout = +1
      10'b0010000110: o_lut = 11'b11011100110;  // D.06.4, RDin = -1, RDout = +1
      10'b0010000111: o_lut = 11'b11011000111;  // D.07.4, RDin = -1, RDout = +1
      10'b0010001000: o_lut = 11'b00100100111;  // D.08.4, RDin = -1, RDout = -1
      10'b0010001001: o_lut = 11'b11011101001;  // D.09.4, RDin = -1, RDout = +1
      10'b0010001010: o_lut = 11'b11011101010;  // D.10.4, RDin = -1, RDout = +1
      10'b0010001011: o_lut = 11'b11011001011;  // D.11.4, RDin = -1, RDout = +1
      10'b0010001100: o_lut = 11'b11011101100;  // D.12.4, RDin = -1, RDout = +1
      10'b0010001101: o_lut = 11'b11011001101;  // D.13.4, RDin = -1, RDout = +1
      10'b0010001110: o_lut = 11'b11011001110;  // D.14.4, RDin = -1, RDout = +1
      10'b0010001111: o_lut = 11'b00100111010;  // D.15.4, RDin = -1, RDout = -1
      10'b0010010000: o_lut = 11'b00100110110;  // D.16.4, RDin = -1, RDout = -1
      10'b0010010001: o_lut = 11'b11011110001;  // D.17.4, RDin = -1, RDout = +1
      10'b0010010010: o_lut = 11'b11011110010;  // D.18.4, RDin = -1, RDout = +1
      10'b0010010011: o_lut = 11'b11011010011;  // D.19.4, RDin = -1, RDout = +1
      10'b0010010100: o_lut = 11'b11011110100;  // D.20.4, RDin = -1, RDout = +1
      10'b0010010101: o_lut = 11'b11011010101;  // D.21.4, RDin = -1, RDout = +1
      10'b0010010110: o_lut = 11'b11011010110;  // D.22.4, RDin = -1, RDout = +1
      10'b0010010111: o_lut = 11'b00100010111;  // D.23.4, RDin = -1, RDout = -1
      10'b0010011000: o_lut = 11'b00100110011;  // D.24.4, RDin = -1, RDout = -1
      10'b0010011001: o_lut = 11'b11011011001;  // D.25.4, RDin = -1, RDout = +1
      10'b0010011010: o_lut = 11'b11011011010;  // D.26.4, RDin = -1, RDout = +1
      10'b0010011011: o_lut = 11'b00100011011;  // D.27.4, RDin = -1, RDout = -1
      10'b0010011100: o_lut = 11'b11011001110;  // D.28.4, RDin = -1, RDout = +1
      10'b0010011101: o_lut = 11'b00100011101;  // D.29.4, RDin = -1, RDout = -1
      10'b0010011110: o_lut = 11'b00100011110;  // D.30.4, RDin = -1, RDout = -1
      10'b0010011111: o_lut = 11'b00100110101;  // D.31.4, RDin = -1, RDout = -1
      10'b0010100000: o_lut = 11'b10101111001;  // D.00.5, RDin = -1, RDout = +1
      10'b0010100001: o_lut = 11'b10101101110;  // D.01.5, RDin = -1, RDout = +1
      10'b0010100010: o_lut = 11'b10101101101;  // D.02.5, RDin = -1, RDout = +1
      10'b0010100011: o_lut = 11'b00101100011;  // D.03.5, RDin = -1, RDout = -1
      10'b0010100100: o_lut = 11'b10101101011;  // D.04.5, RDin = -1, RDout = +1
      10'b0010100101: o_lut = 11'b00101100101;  // D.05.5, RDin = -1, RDout = -1
      10'b0010100110: o_lut = 11'b00101100110;  // D.06.5, RDin = -1, RDout = -1
      10'b0010100111: o_lut = 11'b00101000111;  // D.07.5, RDin = -1, RDout = -1
      10'b0010101000: o_lut = 11'b10101100111;  // D.08.5, RDin = -1, RDout = +1
      10'b0010101001: o_lut = 11'b00101101001;  // D.09.5, RDin = -1, RDout = -1
      10'b0010101010: o_lut = 11'b00101101010;  // D.10.5, RDin = -1, RDout = -1
      10'b0010101011: o_lut = 11'b00101001011;  // D.11.5, RDin = -1, RDout = -1
      10'b0010101100: o_lut = 11'b00101101100;  // D.12.5, RDin = -1, RDout = -1
      10'b0010101101: o_lut = 11'b00101001101;  // D.13.5, RDin = -1, RDout = -1
      10'b0010101110: o_lut = 11'b00101001110;  // D.14.5, RDin = -1, RDout = -1
      10'b0010101111: o_lut = 11'b10101111010;  // D.15.5, RDin = -1, RDout = +1
      10'b0010110000: o_lut = 11'b10101110110;  // D.16.5, RDin = -1, RDout = +1
      10'b0010110001: o_lut = 11'b00101110001;  // D.17.5, RDin = -1, RDout = -1
      10'b0010110010: o_lut = 11'b00101110010;  // D.18.5, RDin = -1, RDout = -1
      10'b0010110011: o_lut = 11'b00101010011;  // D.19.5, RDin = -1, RDout = -1
      10'b0010110100: o_lut = 11'b00101110100;  // D.20.5, RDin = -1, RDout = -1
      10'b0010110101: o_lut = 11'b00101010101;  // D.21.5, RDin = -1, RDout = -1
      10'b0010110110: o_lut = 11'b00101010110;  // D.22.5, RDin = -1, RDout = -1
      10'b0010110111: o_lut = 11'b10101010111;  // D.23.5, RDin = -1, RDout = +1
      10'b0010111000: o_lut = 11'b10101110011;  // D.24.5, RDin = -1, RDout = +1
      10'b0010111001: o_lut = 11'b00101011001;  // D.25.5, RDin = -1, RDout = -1
      10'b0010111010: o_lut = 11'b00101011010;  // D.26.5, RDin = -1, RDout = -1
      10'b0010111011: o_lut = 11'b10101011011;  // D.27.5, RDin = -1, RDout = +1
      10'b0010111100: o_lut = 11'b00101001110;  // D.28.5, RDin = -1, RDout = -1
      10'b0010111101: o_lut = 11'b10101011101;  // D.29.5, RDin = -1, RDout = +1
      10'b0010111110: o_lut = 11'b10101011110;  // D.30.5, RDin = -1, RDout = +1
      10'b0010111111: o_lut = 11'b10101110101;  // D.31.5, RDin = -1, RDout = +1
      10'b0011000000: o_lut = 11'b10110111001;  // D.00.6, RDin = -1, RDout = +1
      10'b0011000001: o_lut = 11'b10110101110;  // D.01.6, RDin = -1, RDout = +1
      10'b0011000010: o_lut = 11'b10110101101;  // D.02.6, RDin = -1, RDout = +1
      10'b0011000011: o_lut = 11'b00110100011;  // D.03.6, RDin = -1, RDout = -1
      10'b0011000100: o_lut = 11'b10110101011;  // D.04.6, RDin = -1, RDout = +1
      10'b0011000101: o_lut = 11'b00110100101;  // D.05.6, RDin = -1, RDout = -1
      10'b0011000110: o_lut = 11'b00110100110;  // D.06.6, RDin = -1, RDout = -1
      10'b0011000111: o_lut = 11'b00110000111;  // D.07.6, RDin = -1, RDout = -1
      10'b0011001000: o_lut = 11'b10110100111;  // D.08.6, RDin = -1, RDout = +1
      10'b0011001001: o_lut = 11'b00110101001;  // D.09.6, RDin = -1, RDout = -1
      10'b0011001010: o_lut = 11'b00110101010;  // D.10.6, RDin = -1, RDout = -1
      10'b0011001011: o_lut = 11'b00110001011;  // D.11.6, RDin = -1, RDout = -1
      10'b0011001100: o_lut = 11'b00110101100;  // D.12.6, RDin = -1, RDout = -1
      10'b0011001101: o_lut = 11'b00110001101;  // D.13.6, RDin = -1, RDout = -1
      10'b0011001110: o_lut = 11'b00110001110;  // D.14.6, RDin = -1, RDout = -1
      10'b0011001111: o_lut = 11'b10110111010;  // D.15.6, RDin = -1, RDout = +1
      10'b0011010000: o_lut = 11'b10110110110;  // D.16.6, RDin = -1, RDout = +1
      10'b0011010001: o_lut = 11'b00110110001;  // D.17.6, RDin = -1, RDout = -1
      10'b0011010010: o_lut = 11'b00110110010;  // D.18.6, RDin = -1, RDout = -1
      10'b0011010011: o_lut = 11'b00110010011;  // D.19.6, RDin = -1, RDout = -1
      10'b0011010100: o_lut = 11'b00110110100;  // D.20.6, RDin = -1, RDout = -1
      10'b0011010101: o_lut = 11'b00110010101;  // D.21.6, RDin = -1, RDout = -1
      10'b0011010110: o_lut = 11'b00110010110;  // D.22.6, RDin = -1, RDout = -1
      10'b0011010111: o_lut = 11'b10110010111;  // D.23.6, RDin = -1, RDout = +1
      10'b0011011000: o_lut = 11'b10110110011;  // D.24.6, RDin = -1, RDout = +1
      10'b0011011001: o_lut = 11'b00110011001;  // D.25.6, RDin = -1, RDout = -1
      10'b0011011010: o_lut = 11'b00110011010;  // D.26.6, RDin = -1, RDout = -1
      10'b0011011011: o_lut = 11'b10110011011;  // D.27.6, RDin = -1, RDout = +1
      10'b0011011100: o_lut = 11'b00110001110;  // D.28.6, RDin = -1, RDout = -1
      10'b0011011101: o_lut = 11'b10110011101;  // D.29.6, RDin = -1, RDout = +1
      10'b0011011110: o_lut = 11'b10110011110;  // D.30.6, RDin = -1, RDout = +1
      10'b0011011111: o_lut = 11'b10110110101;  // D.31.6, RDin = -1, RDout = +1
      10'b0011100000: o_lut = 11'b01000111001;  // D.00.7, RDin = -1, RDout = -1
      10'b0011100001: o_lut = 11'b01000101110;  // D.01.7, RDin = -1, RDout = -1
      10'b0011100010: o_lut = 11'b01000101101;  // D.02.7, RDin = -1, RDout = -1
      10'b0011100011: o_lut = 11'b10111100011;  // D.03.7, RDin = -1, RDout = +1
      10'b0011100100: o_lut = 11'b01000101011;  // D.04.7, RDin = -1, RDout = -1
      10'b0011100101: o_lut = 11'b10111100101;  // D.05.7, RDin = -1, RDout = +1
      10'b0011100110: o_lut = 11'b10111100110;  // D.06.7, RDin = -1, RDout = +1
      10'b0011100111: o_lut = 11'b10111000111;  // D.07.7, RDin = -1, RDout = +1
      10'b0011101000: o_lut = 11'b01000100111;  // D.08.7, RDin = -1, RDout = -1
      10'b0011101001: o_lut = 11'b10111101001;  // D.09.7, RDin = -1, RDout = +1
      10'b0011101010: o_lut = 11'b10111101010;  // D.10.7, RDin = -1, RDout = +1
      10'b0011101011: o_lut = 11'b10111001011;  // D.11.7, RDin = -1, RDout = +1
      10'b0011101100: o_lut = 11'b10111101100;  // D.12.7, RDin = -1, RDout = +1
      10'b0011101101: o_lut = 11'b10111001101;  // D.13.7, RDin = -1, RDout = +1
      10'b0011101110: o_lut = 11'b10111001110;  // D.14.7, RDin = -1, RDout = +1
      10'b0011101111: o_lut = 11'b01000111010;  // D.15.7, RDin = -1, RDout = -1
      10'b0011110000: o_lut = 11'b01000110110;  // D.16.7, RDin = -1, RDout = -1
      10'b0011110001: o_lut = 11'b11110110001;  // D.17.7, RDin = -1, RDout = +1
      10'b0011110010: o_lut = 11'b11110110010;  // D.18.7, RDin = -1, RDout = +1
      10'b0011110011: o_lut = 11'b10111010011;  // D.19.7, RDin = -1, RDout = +1
      10'b0011110100: o_lut = 11'b11110110100;  // D.20.7, RDin = -1, RDout = +1
      10'b0011110101: o_lut = 11'b10111010101;  // D.21.7, RDin = -1, RDout = +1
      10'b0011110110: o_lut = 11'b10111010110;  // D.22.7, RDin = -1, RDout = +1
      10'b0011110111: o_lut = 11'b01000010111;  // D.23.7, RDin = -1, RDout = -1
      10'b0011111000: o_lut = 11'b01000110011;  // D.24.7, RDin = -1, RDout = -1
      10'b0011111001: o_lut = 11'b10111011001;  // D.25.7, RDin = -1, RDout = +1
      10'b0011111010: o_lut = 11'b10111011010;  // D.26.7, RDin = -1, RDout = +1
      10'b0011111011: o_lut = 11'b01000011011;  // D.27.7, RDin = -1, RDout = -1
      10'b0011111100: o_lut = 11'b10111001110;  // D.28.7, RDin = -1, RDout = +1
      10'b0011111101: o_lut = 11'b01000011101;  // D.29.7, RDin = -1, RDout = -1
      10'b0011111110: o_lut = 11'b01000011110;  // D.30.7, RDin = -1, RDout = -1
      10'b0011111111: o_lut = 11'b01000110101;  // D.31.7, RDin = -1, RDout = -1
      10'b0100000000: o_lut = 11'b11101000110;  // D.00.0, RDin = +1, RDout = +1
      10'b0100000001: o_lut = 11'b11101010001;  // D.01.0, RDin = +1, RDout = +1
      10'b0100000010: o_lut = 11'b11101010010;  // D.02.0, RDin = +1, RDout = +1
      10'b0100000011: o_lut = 11'b00010100011;  // D.03.0, RDin = +1, RDout = -1
      10'b0100000100: o_lut = 11'b11101010100;  // D.04.0, RDin = +1, RDout = +1
      10'b0100000101: o_lut = 11'b00010100101;  // D.05.0, RDin = +1, RDout = -1
      10'b0100000110: o_lut = 11'b00010100110;  // D.06.0, RDin = +1, RDout = -1
      10'b0100000111: o_lut = 11'b00010111000;  // D.07.0, RDin = +1, RDout = -1
      10'b0100001000: o_lut = 11'b11101011000;  // D.08.0, RDin = +1, RDout = +1
      10'b0100001001: o_lut = 11'b00010101001;  // D.09.0, RDin = +1, RDout = -1
      10'b0100001010: o_lut = 11'b00010101010;  // D.10.0, RDin = +1, RDout = -1
      10'b0100001011: o_lut = 11'b00010001011;  // D.11.0, RDin = +1, RDout = -1
      10'b0100001100: o_lut = 11'b00010101100;  // D.12.0, RDin = +1, RDout = -1
      10'b0100001101: o_lut = 11'b00010001101;  // D.13.0, RDin = +1, RDout = -1
      10'b0100001110: o_lut = 11'b00010001110;  // D.14.0, RDin = +1, RDout = -1
      10'b0100001111: o_lut = 11'b11101000101;  // D.15.0, RDin = +1, RDout = +1
      10'b0100010000: o_lut = 11'b11101001001;  // D.16.0, RDin = +1, RDout = +1
      10'b0100010001: o_lut = 11'b00010110001;  // D.17.0, RDin = +1, RDout = -1
      10'b0100010010: o_lut = 11'b00010110010;  // D.18.0, RDin = +1, RDout = -1
      10'b0100010011: o_lut = 11'b00010010011;  // D.19.0, RDin = +1, RDout = -1
      10'b0100010100: o_lut = 11'b00010110100;  // D.20.0, RDin = +1, RDout = -1
      10'b0100010101: o_lut = 11'b00010010101;  // D.21.0, RDin = +1, RDout = -1
      10'b0100010110: o_lut = 11'b00010010110;  // D.22.0, RDin = +1, RDout = -1
      10'b0100010111: o_lut = 11'b11101101000;  // D.23.0, RDin = +1, RDout = +1
      10'b0100011000: o_lut = 11'b11101001100;  // D.24.0, RDin = +1, RDout = +1
      10'b0100011001: o_lut = 11'b00010011001;  // D.25.0, RDin = +1, RDout = -1
      10'b0100011010: o_lut = 11'b00010011010;  // D.26.0, RDin = +1, RDout = -1
      10'b0100011011: o_lut = 11'b11101100100;  // D.27.0, RDin = +1, RDout = +1
      10'b0100011100: o_lut = 11'b00010001110;  // D.28.0, RDin = +1, RDout = -1
      10'b0100011101: o_lut = 11'b11101100010;  // D.29.0, RDin = +1, RDout = +1
      10'b0100011110: o_lut = 11'b11101100001;  // D.30.0, RDin = +1, RDout = +1
      10'b0100011111: o_lut = 11'b11101001010;  // D.31.0, RDin = +1, RDout = +1
      10'b0100100000: o_lut = 11'b01001000110;  // D.00.1, RDin = +1, RDout = -1
      10'b0100100001: o_lut = 11'b01001010001;  // D.01.1, RDin = +1, RDout = -1
      10'b0100100010: o_lut = 11'b01001010010;  // D.02.1, RDin = +1, RDout = -1
      10'b0100100011: o_lut = 11'b11001100011;  // D.03.1, RDin = +1, RDout = +1
      10'b0100100100: o_lut = 11'b01001010100;  // D.04.1, RDin = +1, RDout = -1
      10'b0100100101: o_lut = 11'b11001100101;  // D.05.1, RDin = +1, RDout = +1
      10'b0100100110: o_lut = 11'b11001100110;  // D.06.1, RDin = +1, RDout = +1
      10'b0100100111: o_lut = 11'b11001111000;  // D.07.1, RDin = +1, RDout = +1
      10'b0100101000: o_lut = 11'b01001011000;  // D.08.1, RDin = +1, RDout = -1
      10'b0100101001: o_lut = 11'b11001101001;  // D.09.1, RDin = +1, RDout = +1
      10'b0100101010: o_lut = 11'b11001101010;  // D.10.1, RDin = +1, RDout = +1
      10'b0100101011: o_lut = 11'b11001001011;  // D.11.1, RDin = +1, RDout = +1
      10'b0100101100: o_lut = 11'b11001101100;  // D.12.1, RDin = +1, RDout = +1
      10'b0100101101: o_lut = 11'b11001001101;  // D.13.1, RDin = +1, RDout = +1
      10'b0100101110: o_lut = 11'b11001001110;  // D.14.1, RDin = +1, RDout = +1
      10'b0100101111: o_lut = 11'b01001000101;  // D.15.1, RDin = +1, RDout = -1
      10'b0100110000: o_lut = 11'b01001001001;  // D.16.1, RDin = +1, RDout = -1
      10'b0100110001: o_lut = 11'b11001110001;  // D.17.1, RDin = +1, RDout = +1
      10'b0100110010: o_lut = 11'b11001110010;  // D.18.1, RDin = +1, RDout = +1
      10'b0100110011: o_lut = 11'b11001010011;  // D.19.1, RDin = +1, RDout = +1
      10'b0100110100: o_lut = 11'b11001110100;  // D.20.1, RDin = +1, RDout = +1
      10'b0100110101: o_lut = 11'b11001010101;  // D.21.1, RDin = +1, RDout = +1
      10'b0100110110: o_lut = 11'b11001010110;  // D.22.1, RDin = +1, RDout = +1
      10'b0100110111: o_lut = 11'b01001101000;  // D.23.1, RDin = +1, RDout = -1
      10'b0100111000: o_lut = 11'b01001001100;  // D.24.1, RDin = +1, RDout = -1
      10'b0100111001: o_lut = 11'b11001011001;  // D.25.1, RDin = +1, RDout = +1
      10'b0100111010: o_lut = 11'b11001011010;  // D.26.1, RDin = +1, RDout = +1
      10'b0100111011: o_lut = 11'b01001100100;  // D.27.1, RDin = +1, RDout = -1
      10'b0100111100: o_lut = 11'b11001001110;  // D.28.1, RDin = +1, RDout = +1
      10'b0100111101: o_lut = 11'b01001100010;  // D.29.1, RDin = +1, RDout = -1
      10'b0100111110: o_lut = 11'b01001100001;  // D.30.1, RDin = +1, RDout = -1
      10'b0100111111: o_lut = 11'b01001001010;  // D.31.1, RDin = +1, RDout = -1
      10'b0101000000: o_lut = 11'b01010000110;  // D.00.2, RDin = +1, RDout = -1
      10'b0101000001: o_lut = 11'b01010010001;  // D.01.2, RDin = +1, RDout = -1
      10'b0101000010: o_lut = 11'b01010010010;  // D.02.2, RDin = +1, RDout = -1
      10'b0101000011: o_lut = 11'b11010100011;  // D.03.2, RDin = +1, RDout = +1
      10'b0101000100: o_lut = 11'b01010010100;  // D.04.2, RDin = +1, RDout = -1
      10'b0101000101: o_lut = 11'b11010100101;  // D.05.2, RDin = +1, RDout = +1
      10'b0101000110: o_lut = 11'b11010100110;  // D.06.2, RDin = +1, RDout = +1
      10'b0101000111: o_lut = 11'b11010111000;  // D.07.2, RDin = +1, RDout = +1
      10'b0101001000: o_lut = 11'b01010011000;  // D.08.2, RDin = +1, RDout = -1
      10'b0101001001: o_lut = 11'b11010101001;  // D.09.2, RDin = +1, RDout = +1
      10'b0101001010: o_lut = 11'b11010101010;  // D.10.2, RDin = +1, RDout = +1
      10'b0101001011: o_lut = 11'b11010001011;  // D.11.2, RDin = +1, RDout = +1
      10'b0101001100: o_lut = 11'b11010101100;  // D.12.2, RDin = +1, RDout = +1
      10'b0101001101: o_lut = 11'b11010001101;  // D.13.2, RDin = +1, RDout = +1
      10'b0101001110: o_lut = 11'b11010001110;  // D.14.2, RDin = +1, RDout = +1
      10'b0101001111: o_lut = 11'b01010000101;  // D.15.2, RDin = +1, RDout = -1
      10'b0101010000: o_lut = 11'b01010001001;  // D.16.2, RDin = +1, RDout = -1
      10'b0101010001: o_lut = 11'b11010110001;  // D.17.2, RDin = +1, RDout = +1
      10'b0101010010: o_lut = 11'b11010110010;  // D.18.2, RDin = +1, RDout = +1
      10'b0101010011: o_lut = 11'b11010010011;  // D.19.2, RDin = +1, RDout = +1
      10'b0101010100: o_lut = 11'b11010110100;  // D.20.2, RDin = +1, RDout = +1
      10'b0101010101: o_lut = 11'b11010010101;  // D.21.2, RDin = +1, RDout = +1
      10'b0101010110: o_lut = 11'b11010010110;  // D.22.2, RDin = +1, RDout = +1
      10'b0101010111: o_lut = 11'b01010101000;  // D.23.2, RDin = +1, RDout = -1
      10'b0101011000: o_lut = 11'b01010001100;  // D.24.2, RDin = +1, RDout = -1
      10'b0101011001: o_lut = 11'b11010011001;  // D.25.2, RDin = +1, RDout = +1
      10'b0101011010: o_lut = 11'b11010011010;  // D.26.2, RDin = +1, RDout = +1
      10'b0101011011: o_lut = 11'b01010100100;  // D.27.2, RDin = +1, RDout = -1
      10'b0101011100: o_lut = 11'b11010001110;  // D.28.2, RDin = +1, RDout = +1
      10'b0101011101: o_lut = 11'b01010100010;  // D.29.2, RDin = +1, RDout = -1
      10'b0101011110: o_lut = 11'b01010100001;  // D.30.2, RDin = +1, RDout = -1
      10'b0101011111: o_lut = 11'b01010001010;  // D.31.2, RDin = +1, RDout = -1
      10'b0101100000: o_lut = 11'b00011000110;  // D.00.3, RDin = +1, RDout = -1
      10'b0101100001: o_lut = 11'b00011010001;  // D.01.3, RDin = +1, RDout = -1
      10'b0101100010: o_lut = 11'b00011010010;  // D.02.3, RDin = +1, RDout = -1
      10'b0101100011: o_lut = 11'b11100100011;  // D.03.3, RDin = +1, RDout = +1
      10'b0101100100: o_lut = 11'b00011010100;  // D.04.3, RDin = +1, RDout = -1
      10'b0101100101: o_lut = 11'b11100100101;  // D.05.3, RDin = +1, RDout = +1
      10'b0101100110: o_lut = 11'b11100100110;  // D.06.3, RDin = +1, RDout = +1
      10'b0101100111: o_lut = 11'b11100111000;  // D.07.3, RDin = +1, RDout = +1
      10'b0101101000: o_lut = 11'b00011011000;  // D.08.3, RDin = +1, RDout = -1
      10'b0101101001: o_lut = 11'b11100101001;  // D.09.3, RDin = +1, RDout = +1
      10'b0101101010: o_lut = 11'b11100101010;  // D.10.3, RDin = +1, RDout = +1
      10'b0101101011: o_lut = 11'b11100001011;  // D.11.3, RDin = +1, RDout = +1
      10'b0101101100: o_lut = 11'b11100101100;  // D.12.3, RDin = +1, RDout = +1
      10'b0101101101: o_lut = 11'b11100001101;  // D.13.3, RDin = +1, RDout = +1
      10'b0101101110: o_lut = 11'b11100001110;  // D.14.3, RDin = +1, RDout = +1
      10'b0101101111: o_lut = 11'b00011000101;  // D.15.3, RDin = +1, RDout = -1
      10'b0101110000: o_lut = 11'b00011001001;  // D.16.3, RDin = +1, RDout = -1
      10'b0101110001: o_lut = 11'b11100110001;  // D.17.3, RDin = +1, RDout = +1
      10'b0101110010: o_lut = 11'b11100110010;  // D.18.3, RDin = +1, RDout = +1
      10'b0101110011: o_lut = 11'b11100010011;  // D.19.3, RDin = +1, RDout = +1
      10'b0101110100: o_lut = 11'b11100110100;  // D.20.3, RDin = +1, RDout = +1
      10'b0101110101: o_lut = 11'b11100010101;  // D.21.3, RDin = +1, RDout = +1
      10'b0101110110: o_lut = 11'b11100010110;  // D.22.3, RDin = +1, RDout = +1
      10'b0101110111: o_lut = 11'b00011101000;  // D.23.3, RDin = +1, RDout = -1
      10'b0101111000: o_lut = 11'b00011001100;  // D.24.3, RDin = +1, RDout = -1
      10'b0101111001: o_lut = 11'b11100011001;  // D.25.3, RDin = +1, RDout = +1
      10'b0101111010: o_lut = 11'b11100011010;  // D.26.3, RDin = +1, RDout = +1
      10'b0101111011: o_lut = 11'b00011100100;  // D.27.3, RDin = +1, RDout = -1
      10'b0101111100: o_lut = 11'b11100001110;  // D.28.3, RDin = +1, RDout = +1
      10'b0101111101: o_lut = 11'b00011100010;  // D.29.3, RDin = +1, RDout = -1
      10'b0101111110: o_lut = 11'b00011100001;  // D.30.3, RDin = +1, RDout = -1
      10'b0101111111: o_lut = 11'b00011001010;  // D.31.3, RDin = +1, RDout = -1
      10'b0110000000: o_lut = 11'b11011000110;  // D.00.4, RDin = +1, RDout = +1
      10'b0110000001: o_lut = 11'b11011010001;  // D.01.4, RDin = +1, RDout = +1
      10'b0110000010: o_lut = 11'b11011010010;  // D.02.4, RDin = +1, RDout = +1
      10'b0110000011: o_lut = 11'b00100100011;  // D.03.4, RDin = +1, RDout = -1
      10'b0110000100: o_lut = 11'b11011010100;  // D.04.4, RDin = +1, RDout = +1
      10'b0110000101: o_lut = 11'b00100100101;  // D.05.4, RDin = +1, RDout = -1
      10'b0110000110: o_lut = 11'b00100100110;  // D.06.4, RDin = +1, RDout = -1
      10'b0110000111: o_lut = 11'b00100111000;  // D.07.4, RDin = +1, RDout = -1
      10'b0110001000: o_lut = 11'b11011011000;  // D.08.4, RDin = +1, RDout = +1
      10'b0110001001: o_lut = 11'b00100101001;  // D.09.4, RDin = +1, RDout = -1
      10'b0110001010: o_lut = 11'b00100101010;  // D.10.4, RDin = +1, RDout = -1
      10'b0110001011: o_lut = 11'b00100001011;  // D.11.4, RDin = +1, RDout = -1
      10'b0110001100: o_lut = 11'b00100101100;  // D.12.4, RDin = +1, RDout = -1
      10'b0110001101: o_lut = 11'b00100001101;  // D.13.4, RDin = +1, RDout = -1
      10'b0110001110: o_lut = 11'b00100001110;  // D.14.4, RDin = +1, RDout = -1
      10'b0110001111: o_lut = 11'b11011000101;  // D.15.4, RDin = +1, RDout = +1
      10'b0110010000: o_lut = 11'b11011001001;  // D.16.4, RDin = +1, RDout = +1
      10'b0110010001: o_lut = 11'b00100110001;  // D.17.4, RDin = +1, RDout = -1
      10'b0110010010: o_lut = 11'b00100110010;  // D.18.4, RDin = +1, RDout = -1
      10'b0110010011: o_lut = 11'b00100010011;  // D.19.4, RDin = +1, RDout = -1
      10'b0110010100: o_lut = 11'b00100110100;  // D.20.4, RDin = +1, RDout = -1
      10'b0110010101: o_lut = 11'b00100010101;  // D.21.4, RDin = +1, RDout = -1
      10'b0110010110: o_lut = 11'b00100010110;  // D.22.4, RDin = +1, RDout = -1
      10'b0110010111: o_lut = 11'b11011101000;  // D.23.4, RDin = +1, RDout = +1
      10'b0110011000: o_lut = 11'b11011001100;  // D.24.4, RDin = +1, RDout = +1
      10'b0110011001: o_lut = 11'b00100011001;  // D.25.4, RDin = +1, RDout = -1
      10'b0110011010: o_lut = 11'b00100011010;  // D.26.4, RDin = +1, RDout = -1
      10'b0110011011: o_lut = 11'b11011100100;  // D.27.4, RDin = +1, RDout = +1
      10'b0110011100: o_lut = 11'b00100001110;  // D.28.4, RDin = +1, RDout = -1
      10'b0110011101: o_lut = 11'b11011100010;  // D.29.4, RDin = +1, RDout = +1
      10'b0110011110: o_lut = 11'b11011100001;  // D.30.4, RDin = +1, RDout = +1
      10'b0110011111: o_lut = 11'b11011001010;  // D.31.4, RDin = +1, RDout = +1
      10'b0110100000: o_lut = 11'b00101000110;  // D.00.5, RDin = +1, RDout = -1
      10'b0110100001: o_lut = 11'b00101010001;  // D.01.5, RDin = +1, RDout = -1
      10'b0110100010: o_lut = 11'b00101010010;  // D.02.5, RDin = +1, RDout = -1
      10'b0110100011: o_lut = 11'b10101100011;  // D.03.5, RDin = +1, RDout = +1
      10'b0110100100: o_lut = 11'b00101010100;  // D.04.5, RDin = +1, RDout = -1
      10'b0110100101: o_lut = 11'b10101100101;  // D.05.5, RDin = +1, RDout = +1
      10'b0110100110: o_lut = 11'b10101100110;  // D.06.5, RDin = +1, RDout = +1
      10'b0110100111: o_lut = 11'b10101111000;  // D.07.5, RDin = +1, RDout = +1
      10'b0110101000: o_lut = 11'b00101011000;  // D.08.5, RDin = +1, RDout = -1
      10'b0110101001: o_lut = 11'b10101101001;  // D.09.5, RDin = +1, RDout = +1
      10'b0110101010: o_lut = 11'b10101101010;  // D.10.5, RDin = +1, RDout = +1
      10'b0110101011: o_lut = 11'b10101001011;  // D.11.5, RDin = +1, RDout = +1
      10'b0110101100: o_lut = 11'b10101101100;  // D.12.5, RDin = +1, RDout = +1
      10'b0110101101: o_lut = 11'b10101001101;  // D.13.5, RDin = +1, RDout = +1
      10'b0110101110: o_lut = 11'b10101001110;  // D.14.5, RDin = +1, RDout = +1
      10'b0110101111: o_lut = 11'b00101000101;  // D.15.5, RDin = +1, RDout = -1
      10'b0110110000: o_lut = 11'b00101001001;  // D.16.5, RDin = +1, RDout = -1
      10'b0110110001: o_lut = 11'b10101110001;  // D.17.5, RDin = +1, RDout = +1
      10'b0110110010: o_lut = 11'b10101110010;  // D.18.5, RDin = +1, RDout = +1
      10'b0110110011: o_lut = 11'b10101010011;  // D.19.5, RDin = +1, RDout = +1
      10'b0110110100: o_lut = 11'b10101110100;  // D.20.5, RDin = +1, RDout = +1
      10'b0110110101: o_lut = 11'b10101010101;  // D.21.5, RDin = +1, RDout = +1
      10'b0110110110: o_lut = 11'b10101010110;  // D.22.5, RDin = +1, RDout = +1
      10'b0110110111: o_lut = 11'b00101101000;  // D.23.5, RDin = +1, RDout = -1
      10'b0110111000: o_lut = 11'b00101001100;  // D.24.5, RDin = +1, RDout = -1
      10'b0110111001: o_lut = 11'b10101011001;  // D.25.5, RDin = +1, RDout = +1
      10'b0110111010: o_lut = 11'b10101011010;  // D.26.5, RDin = +1, RDout = +1
      10'b0110111011: o_lut = 11'b00101100100;  // D.27.5, RDin = +1, RDout = -1
      10'b0110111100: o_lut = 11'b10101001110;  // D.28.5, RDin = +1, RDout = +1
      10'b0110111101: o_lut = 11'b00101100010;  // D.29.5, RDin = +1, RDout = -1
      10'b0110111110: o_lut = 11'b00101100001;  // D.30.5, RDin = +1, RDout = -1
      10'b0110111111: o_lut = 11'b00101001010;  // D.31.5, RDin = +1, RDout = -1
      10'b0111000000: o_lut = 11'b00110000110;  // D.00.6, RDin = +1, RDout = -1
      10'b0111000001: o_lut = 11'b00110010001;  // D.01.6, RDin = +1, RDout = -1
      10'b0111000010: o_lut = 11'b00110010010;  // D.02.6, RDin = +1, RDout = -1
      10'b0111000011: o_lut = 11'b10110100011;  // D.03.6, RDin = +1, RDout = +1
      10'b0111000100: o_lut = 11'b00110010100;  // D.04.6, RDin = +1, RDout = -1
      10'b0111000101: o_lut = 11'b10110100101;  // D.05.6, RDin = +1, RDout = +1
      10'b0111000110: o_lut = 11'b10110100110;  // D.06.6, RDin = +1, RDout = +1
      10'b0111000111: o_lut = 11'b10110111000;  // D.07.6, RDin = +1, RDout = +1
      10'b0111001000: o_lut = 11'b00110011000;  // D.08.6, RDin = +1, RDout = -1
      10'b0111001001: o_lut = 11'b10110101001;  // D.09.6, RDin = +1, RDout = +1
      10'b0111001010: o_lut = 11'b10110101010;  // D.10.6, RDin = +1, RDout = +1
      10'b0111001011: o_lut = 11'b10110001011;  // D.11.6, RDin = +1, RDout = +1
      10'b0111001100: o_lut = 11'b10110101100;  // D.12.6, RDin = +1, RDout = +1
      10'b0111001101: o_lut = 11'b10110001101;  // D.13.6, RDin = +1, RDout = +1
      10'b0111001110: o_lut = 11'b10110001110;  // D.14.6, RDin = +1, RDout = +1
      10'b0111001111: o_lut = 11'b00110000101;  // D.15.6, RDin = +1, RDout = -1
      10'b0111010000: o_lut = 11'b00110001001;  // D.16.6, RDin = +1, RDout = -1
      10'b0111010001: o_lut = 11'b10110110001;  // D.17.6, RDin = +1, RDout = +1
      10'b0111010010: o_lut = 11'b10110110010;  // D.18.6, RDin = +1, RDout = +1
      10'b0111010011: o_lut = 11'b10110010011;  // D.19.6, RDin = +1, RDout = +1
      10'b0111010100: o_lut = 11'b10110110100;  // D.20.6, RDin = +1, RDout = +1
      10'b0111010101: o_lut = 11'b10110010101;  // D.21.6, RDin = +1, RDout = +1
      10'b0111010110: o_lut = 11'b10110010110;  // D.22.6, RDin = +1, RDout = +1
      10'b0111010111: o_lut = 11'b00110101000;  // D.23.6, RDin = +1, RDout = -1
      10'b0111011000: o_lut = 11'b00110001100;  // D.24.6, RDin = +1, RDout = -1
      10'b0111011001: o_lut = 11'b10110011001;  // D.25.6, RDin = +1, RDout = +1
      10'b0111011010: o_lut = 11'b10110011010;  // D.26.6, RDin = +1, RDout = +1
      10'b0111011011: o_lut = 11'b00110100100;  // D.27.6, RDin = +1, RDout = -1
      10'b0111011100: o_lut = 11'b10110001110;  // D.28.6, RDin = +1, RDout = +1
      10'b0111011101: o_lut = 11'b00110100010;  // D.29.6, RDin = +1, RDout = -1
      10'b0111011110: o_lut = 11'b00110100001;  // D.30.6, RDin = +1, RDout = -1
      10'b0111011111: o_lut = 11'b00110001010;  // D.31.6, RDin = +1, RDout = -1
      10'b0111100000: o_lut = 11'b10111000110;  // D.00.7, RDin = +1, RDout = +1
      10'b0111100001: o_lut = 11'b10111010001;  // D.01.7, RDin = +1, RDout = +1
      10'b0111100010: o_lut = 11'b10111010010;  // D.02.7, RDin = +1, RDout = +1
      10'b0111100011: o_lut = 11'b01000100011;  // D.03.7, RDin = +1, RDout = -1
      10'b0111100100: o_lut = 11'b10111010100;  // D.04.7, RDin = +1, RDout = +1
      10'b0111100101: o_lut = 11'b01000100101;  // D.05.7, RDin = +1, RDout = -1
      10'b0111100110: o_lut = 11'b01000100110;  // D.06.7, RDin = +1, RDout = -1
      10'b0111100111: o_lut = 11'b01000111000;  // D.07.7, RDin = +1, RDout = -1
      10'b0111101000: o_lut = 11'b10111011000;  // D.08.7, RDin = +1, RDout = +1
      10'b0111101001: o_lut = 11'b01000101001;  // D.09.7, RDin = +1, RDout = -1
      10'b0111101010: o_lut = 11'b01000101010;  // D.10.7, RDin = +1, RDout = -1
      10'b0111101011: o_lut = 11'b00001001011;  // D.11.7, RDin = +1, RDout = -1
      10'b0111101100: o_lut = 11'b01000101100;  // D.12.7, RDin = +1, RDout = -1
      10'b0111101101: o_lut = 11'b00001001101;  // D.13.7, RDin = +1, RDout = -1
      10'b0111101110: o_lut = 11'b00001001110;  // D.14.7, RDin = +1, RDout = -1
      10'b0111101111: o_lut = 11'b10111000101;  // D.15.7, RDin = +1, RDout = +1
      10'b0111110000: o_lut = 11'b10111001001;  // D.16.7, RDin = +1, RDout = +1
      10'b0111110001: o_lut = 11'b01000110001;  // D.17.7, RDin = +1, RDout = -1
      10'b0111110010: o_lut = 11'b01000110010;  // D.18.7, RDin = +1, RDout = -1
      10'b0111110011: o_lut = 11'b01000010011;  // D.19.7, RDin = +1, RDout = -1
      10'b0111110100: o_lut = 11'b01000110100;  // D.20.7, RDin = +1, RDout = -1
      10'b0111110101: o_lut = 11'b01000010101;  // D.21.7, RDin = +1, RDout = -1
      10'b0111110110: o_lut = 11'b01000010110;  // D.22.7, RDin = +1, RDout = -1
      10'b0111110111: o_lut = 11'b10111101000;  // D.23.7, RDin = +1, RDout = +1
      10'b0111111000: o_lut = 11'b10111001100;  // D.24.7, RDin = +1, RDout = +1
      10'b0111111001: o_lut = 11'b01000011001;  // D.25.7, RDin = +1, RDout = -1
      10'b0111111010: o_lut = 11'b01000011010;  // D.26.7, RDin = +1, RDout = -1
      10'b0111111011: o_lut = 11'b10111100100;  // D.27.7, RDin = +1, RDout = +1
      10'b0111111100: o_lut = 11'b01000001110;  // D.28.7, RDin = +1, RDout = -1
      10'b0111111101: o_lut = 11'b10111100010;  // D.29.7, RDin = +1, RDout = +1
      10'b0111111110: o_lut = 11'b10111100001;  // D.30.7, RDin = +1, RDout = +1
      10'b0111111111: o_lut = 11'b10111001010;  // D.31.7, RDin = +1, RDout = +1
      10'b1000000000: o_lut = 11'b00010111001;  // K.00.0, RDin = -1, RDout = -1
      10'b1000000001: o_lut = 11'b00010101110;  // K.01.0, RDin = -1, RDout = -1
      10'b1000000010: o_lut = 11'b00010101101;  // K.02.0, RDin = -1, RDout = -1
      10'b1000000011: o_lut = 11'b11101100011;  // K.03.0, RDin = -1, RDout = +1
      10'b1000000100: o_lut = 11'b00010101011;  // K.04.0, RDin = -1, RDout = -1
      10'b1000000101: o_lut = 11'b11101100101;  // K.05.0, RDin = -1, RDout = +1
      10'b1000000110: o_lut = 11'b11101100110;  // K.06.0, RDin = -1, RDout = +1
      10'b1000000111: o_lut = 11'b11101000111;  // K.07.0, RDin = -1, RDout = +1
      10'b1000001000: o_lut = 11'b00010100111;  // K.08.0, RDin = -1, RDout = -1
      10'b1000001001: o_lut = 11'b11101101001;  // K.09.0, RDin = -1, RDout = +1
      10'b1000001010: o_lut = 11'b11101101010;  // K.10.0, RDin = -1, RDout = +1
      10'b1000001011: o_lut = 11'b11101001011;  // K.11.0, RDin = -1, RDout = +1
      10'b1000001100: o_lut = 11'b11101101100;  // K.12.0, RDin = -1, RDout = +1
      10'b1000001101: o_lut = 11'b11101001101;  // K.13.0, RDin = -1, RDout = +1
      10'b1000001110: o_lut = 11'b11101001110;  // K.14.0, RDin = -1, RDout = +1
      10'b1000001111: o_lut = 11'b00010111010;  // K.15.0, RDin = -1, RDout = -1
      10'b1000010000: o_lut = 11'b00010110110;  // K.16.0, RDin = -1, RDout = -1
      10'b1000010001: o_lut = 11'b11101110001;  // K.17.0, RDin = -1, RDout = +1
      10'b1000010010: o_lut = 11'b11101110010;  // K.18.0, RDin = -1, RDout = +1
      10'b1000010011: o_lut = 11'b11101010011;  // K.19.0, RDin = -1, RDout = +1
      10'b1000010100: o_lut = 11'b11101110100;  // K.20.0, RDin = -1, RDout = +1
      10'b1000010101: o_lut = 11'b11101010101;  // K.21.0, RDin = -1, RDout = +1
      10'b1000010110: o_lut = 11'b11101010110;  // K.22.0, RDin = -1, RDout = +1
      10'b1000010111: o_lut = 11'b00010010111;  // K.23.0, RDin = -1, RDout = -1
      10'b1000011000: o_lut = 11'b00010110011;  // K.24.0, RDin = -1, RDout = -1
      10'b1000011001: o_lut = 11'b11101011001;  // K.25.0, RDin = -1, RDout = +1
      10'b1000011010: o_lut = 11'b11101011010;  // K.26.0, RDin = -1, RDout = +1
      10'b1000011011: o_lut = 11'b00010011011;  // K.27.0, RDin = -1, RDout = -1
      10'b1000011100: o_lut = 11'b00010111100;  // K.28.0, RDin = -1, RDout = -1
      10'b1000011101: o_lut = 11'b00010011101;  // K.29.0, RDin = -1, RDout = -1
      10'b1000011110: o_lut = 11'b00010011110;  // K.30.0, RDin = -1, RDout = -1
      10'b1000011111: o_lut = 11'b00010110101;  // K.31.0, RDin = -1, RDout = -1
      10'b1000100000: o_lut = 11'b11001111001;  // K.00.1, RDin = -1, RDout = +1
      10'b1000100001: o_lut = 11'b11001101110;  // K.01.1, RDin = -1, RDout = +1
      10'b1000100010: o_lut = 11'b11001101101;  // K.02.1, RDin = -1, RDout = +1
      10'b1000100011: o_lut = 11'b00110100011;  // K.03.1, RDin = -1, RDout = -1
      10'b1000100100: o_lut = 11'b11001101011;  // K.04.1, RDin = -1, RDout = +1
      10'b1000100101: o_lut = 11'b00110100101;  // K.05.1, RDin = -1, RDout = -1
      10'b1000100110: o_lut = 11'b00110100110;  // K.06.1, RDin = -1, RDout = -1
      10'b1000100111: o_lut = 11'b00110000111;  // K.07.1, RDin = -1, RDout = -1
      10'b1000101000: o_lut = 11'b11001100111;  // K.08.1, RDin = -1, RDout = +1
      10'b1000101001: o_lut = 11'b00110101001;  // K.09.1, RDin = -1, RDout = -1
      10'b1000101010: o_lut = 11'b00110101010;  // K.10.1, RDin = -1, RDout = -1
      10'b1000101011: o_lut = 11'b00110001011;  // K.11.1, RDin = -1, RDout = -1
      10'b1000101100: o_lut = 11'b00110101100;  // K.12.1, RDin = -1, RDout = -1
      10'b1000101101: o_lut = 11'b00110001101;  // K.13.1, RDin = -1, RDout = -1
      10'b1000101110: o_lut = 11'b00110001110;  // K.14.1, RDin = -1, RDout = -1
      10'b1000101111: o_lut = 11'b11001111010;  // K.15.1, RDin = -1, RDout = +1
      10'b1000110000: o_lut = 11'b11001110110;  // K.16.1, RDin = -1, RDout = +1
      10'b1000110001: o_lut = 11'b00110110001;  // K.17.1, RDin = -1, RDout = -1
      10'b1000110010: o_lut = 11'b00110110010;  // K.18.1, RDin = -1, RDout = -1
      10'b1000110011: o_lut = 11'b00110010011;  // K.19.1, RDin = -1, RDout = -1
      10'b1000110100: o_lut = 11'b00110110100;  // K.20.1, RDin = -1, RDout = -1
      10'b1000110101: o_lut = 11'b00110010101;  // K.21.1, RDin = -1, RDout = -1
      10'b1000110110: o_lut = 11'b00110010110;  // K.22.1, RDin = -1, RDout = -1
      10'b1000110111: o_lut = 11'b11001010111;  // K.23.1, RDin = -1, RDout = +1
      10'b1000111000: o_lut = 11'b11001110011;  // K.24.1, RDin = -1, RDout = +1
      10'b1000111001: o_lut = 11'b00110011001;  // K.25.1, RDin = -1, RDout = -1
      10'b1000111010: o_lut = 11'b00110011010;  // K.26.1, RDin = -1, RDout = -1
      10'b1000111011: o_lut = 11'b11001011011;  // K.27.1, RDin = -1, RDout = +1
      10'b1000111100: o_lut = 11'b11001111100;  // K.28.1, RDin = -1, RDout = +1
      10'b1000111101: o_lut = 11'b11001011101;  // K.29.1, RDin = -1, RDout = +1
      10'b1000111110: o_lut = 11'b11001011110;  // K.30.1, RDin = -1, RDout = +1
      10'b1000111111: o_lut = 11'b11001110101;  // K.31.1, RDin = -1, RDout = +1
      10'b1001000000: o_lut = 11'b11010111001;  // K.00.2, RDin = -1, RDout = +1
      10'b1001000001: o_lut = 11'b11010101110;  // K.01.2, RDin = -1, RDout = +1
      10'b1001000010: o_lut = 11'b11010101101;  // K.02.2, RDin = -1, RDout = +1
      10'b1001000011: o_lut = 11'b00101100011;  // K.03.2, RDin = -1, RDout = -1
      10'b1001000100: o_lut = 11'b11010101011;  // K.04.2, RDin = -1, RDout = +1
      10'b1001000101: o_lut = 11'b00101100101;  // K.05.2, RDin = -1, RDout = -1
      10'b1001000110: o_lut = 11'b00101100110;  // K.06.2, RDin = -1, RDout = -1
      10'b1001000111: o_lut = 11'b00101000111;  // K.07.2, RDin = -1, RDout = -1
      10'b1001001000: o_lut = 11'b11010100111;  // K.08.2, RDin = -1, RDout = +1
      10'b1001001001: o_lut = 11'b00101101001;  // K.09.2, RDin = -1, RDout = -1
      10'b1001001010: o_lut = 11'b00101101010;  // K.10.2, RDin = -1, RDout = -1
      10'b1001001011: o_lut = 11'b00101001011;  // K.11.2, RDin = -1, RDout = -1
      10'b1001001100: o_lut = 11'b00101101100;  // K.12.2, RDin = -1, RDout = -1
      10'b1001001101: o_lut = 11'b00101001101;  // K.13.2, RDin = -1, RDout = -1
      10'b1001001110: o_lut = 11'b00101001110;  // K.14.2, RDin = -1, RDout = -1
      10'b1001001111: o_lut = 11'b11010111010;  // K.15.2, RDin = -1, RDout = +1
      10'b1001010000: o_lut = 11'b11010110110;  // K.16.2, RDin = -1, RDout = +1
      10'b1001010001: o_lut = 11'b00101110001;  // K.17.2, RDin = -1, RDout = -1
      10'b1001010010: o_lut = 11'b00101110010;  // K.18.2, RDin = -1, RDout = -1
      10'b1001010011: o_lut = 11'b00101010011;  // K.19.2, RDin = -1, RDout = -1
      10'b1001010100: o_lut = 11'b00101110100;  // K.20.2, RDin = -1, RDout = -1
      10'b1001010101: o_lut = 11'b00101010101;  // K.21.2, RDin = -1, RDout = -1
      10'b1001010110: o_lut = 11'b00101010110;  // K.22.2, RDin = -1, RDout = -1
      10'b1001010111: o_lut = 11'b11010010111;  // K.23.2, RDin = -1, RDout = +1
      10'b1001011000: o_lut = 11'b11010110011;  // K.24.2, RDin = -1, RDout = +1
      10'b1001011001: o_lut = 11'b00101011001;  // K.25.2, RDin = -1, RDout = -1
      10'b1001011010: o_lut = 11'b00101011010;  // K.26.2, RDin = -1, RDout = -1
      10'b1001011011: o_lut = 11'b11010011011;  // K.27.2, RDin = -1, RDout = +1
      10'b1001011100: o_lut = 11'b11010111100;  // K.28.2, RDin = -1, RDout = +1
      10'b1001011101: o_lut = 11'b11010011101;  // K.29.2, RDin = -1, RDout = +1
      10'b1001011110: o_lut = 11'b11010011110;  // K.30.2, RDin = -1, RDout = +1
      10'b1001011111: o_lut = 11'b11010110101;  // K.31.2, RDin = -1, RDout = +1
      10'b1001100000: o_lut = 11'b11100111001;  // K.00.3, RDin = -1, RDout = +1
      10'b1001100001: o_lut = 11'b11100101110;  // K.01.3, RDin = -1, RDout = +1
      10'b1001100010: o_lut = 11'b11100101101;  // K.02.3, RDin = -1, RDout = +1
      10'b1001100011: o_lut = 11'b00011100011;  // K.03.3, RDin = -1, RDout = -1
      10'b1001100100: o_lut = 11'b11100101011;  // K.04.3, RDin = -1, RDout = +1
      10'b1001100101: o_lut = 11'b00011100101;  // K.05.3, RDin = -1, RDout = -1
      10'b1001100110: o_lut = 11'b00011100110;  // K.06.3, RDin = -1, RDout = -1
      10'b1001100111: o_lut = 11'b00011000111;  // K.07.3, RDin = -1, RDout = -1
      10'b1001101000: o_lut = 11'b11100100111;  // K.08.3, RDin = -1, RDout = +1
      10'b1001101001: o_lut = 11'b00011101001;  // K.09.3, RDin = -1, RDout = -1
      10'b1001101010: o_lut = 11'b00011101010;  // K.10.3, RDin = -1, RDout = -1
      10'b1001101011: o_lut = 11'b00011001011;  // K.11.3, RDin = -1, RDout = -1
      10'b1001101100: o_lut = 11'b00011101100;  // K.12.3, RDin = -1, RDout = -1
      10'b1001101101: o_lut = 11'b00011001101;  // K.13.3, RDin = -1, RDout = -1
      10'b1001101110: o_lut = 11'b00011001110;  // K.14.3, RDin = -1, RDout = -1
      10'b1001101111: o_lut = 11'b11100111010;  // K.15.3, RDin = -1, RDout = +1
      10'b1001110000: o_lut = 11'b11100110110;  // K.16.3, RDin = -1, RDout = +1
      10'b1001110001: o_lut = 11'b00011110001;  // K.17.3, RDin = -1, RDout = -1
      10'b1001110010: o_lut = 11'b00011110010;  // K.18.3, RDin = -1, RDout = -1
      10'b1001110011: o_lut = 11'b00011010011;  // K.19.3, RDin = -1, RDout = -1
      10'b1001110100: o_lut = 11'b00011110100;  // K.20.3, RDin = -1, RDout = -1
      10'b1001110101: o_lut = 11'b00011010101;  // K.21.3, RDin = -1, RDout = -1
      10'b1001110110: o_lut = 11'b00011010110;  // K.22.3, RDin = -1, RDout = -1
      10'b1001110111: o_lut = 11'b11100010111;  // K.23.3, RDin = -1, RDout = +1
      10'b1001111000: o_lut = 11'b11100110011;  // K.24.3, RDin = -1, RDout = +1
      10'b1001111001: o_lut = 11'b00011011001;  // K.25.3, RDin = -1, RDout = -1
      10'b1001111010: o_lut = 11'b00011011010;  // K.26.3, RDin = -1, RDout = -1
      10'b1001111011: o_lut = 11'b11100011011;  // K.27.3, RDin = -1, RDout = +1
      10'b1001111100: o_lut = 11'b11100111100;  // K.28.3, RDin = -1, RDout = +1
      10'b1001111101: o_lut = 11'b11100011101;  // K.29.3, RDin = -1, RDout = +1
      10'b1001111110: o_lut = 11'b11100011110;  // K.30.3, RDin = -1, RDout = +1
      10'b1001111111: o_lut = 11'b11100110101;  // K.31.3, RDin = -1, RDout = +1
      10'b1010000000: o_lut = 11'b00100111001;  // K.00.4, RDin = -1, RDout = -1
      10'b1010000001: o_lut = 11'b00100101110;  // K.01.4, RDin = -1, RDout = -1
      10'b1010000010: o_lut = 11'b00100101101;  // K.02.4, RDin = -1, RDout = -1
      10'b1010000011: o_lut = 11'b11011100011;  // K.03.4, RDin = -1, RDout = +1
      10'b1010000100: o_lut = 11'b00100101011;  // K.04.4, RDin = -1, RDout = -1
      10'b1010000101: o_lut = 11'b11011100101;  // K.05.4, RDin = -1, RDout = +1
      10'b1010000110: o_lut = 11'b11011100110;  // K.06.4, RDin = -1, RDout = +1
      10'b1010000111: o_lut = 11'b11011000111;  // K.07.4, RDin = -1, RDout = +1
      10'b1010001000: o_lut = 11'b00100100111;  // K.08.4, RDin = -1, RDout = -1
      10'b1010001001: o_lut = 11'b11011101001;  // K.09.4, RDin = -1, RDout = +1
      10'b1010001010: o_lut = 11'b11011101010;  // K.10.4, RDin = -1, RDout = +1
      10'b1010001011: o_lut = 11'b11011001011;  // K.11.4, RDin = -1, RDout = +1
      10'b1010001100: o_lut = 11'b11011101100;  // K.12.4, RDin = -1, RDout = +1
      10'b1010001101: o_lut = 11'b11011001101;  // K.13.4, RDin = -1, RDout = +1
      10'b1010001110: o_lut = 11'b11011001110;  // K.14.4, RDin = -1, RDout = +1
      10'b1010001111: o_lut = 11'b00100111010;  // K.15.4, RDin = -1, RDout = -1
      10'b1010010000: o_lut = 11'b00100110110;  // K.16.4, RDin = -1, RDout = -1
      10'b1010010001: o_lut = 11'b11011110001;  // K.17.4, RDin = -1, RDout = +1
      10'b1010010010: o_lut = 11'b11011110010;  // K.18.4, RDin = -1, RDout = +1
      10'b1010010011: o_lut = 11'b11011010011;  // K.19.4, RDin = -1, RDout = +1
      10'b1010010100: o_lut = 11'b11011110100;  // K.20.4, RDin = -1, RDout = +1
      10'b1010010101: o_lut = 11'b11011010101;  // K.21.4, RDin = -1, RDout = +1
      10'b1010010110: o_lut = 11'b11011010110;  // K.22.4, RDin = -1, RDout = +1
      10'b1010010111: o_lut = 11'b00100010111;  // K.23.4, RDin = -1, RDout = -1
      10'b1010011000: o_lut = 11'b00100110011;  // K.24.4, RDin = -1, RDout = -1
      10'b1010011001: o_lut = 11'b11011011001;  // K.25.4, RDin = -1, RDout = +1
      10'b1010011010: o_lut = 11'b11011011010;  // K.26.4, RDin = -1, RDout = +1
      10'b1010011011: o_lut = 11'b00100011011;  // K.27.4, RDin = -1, RDout = -1
      10'b1010011100: o_lut = 11'b00100111100;  // K.28.4, RDin = -1, RDout = -1
      10'b1010011101: o_lut = 11'b00100011101;  // K.29.4, RDin = -1, RDout = -1
      10'b1010011110: o_lut = 11'b00100011110;  // K.30.4, RDin = -1, RDout = -1
      10'b1010011111: o_lut = 11'b00100110101;  // K.31.4, RDin = -1, RDout = -1
      10'b1010100000: o_lut = 11'b10101111001;  // K.00.5, RDin = -1, RDout = +1
      10'b1010100001: o_lut = 11'b10101101110;  // K.01.5, RDin = -1, RDout = +1
      10'b1010100010: o_lut = 11'b10101101101;  // K.02.5, RDin = -1, RDout = +1
      10'b1010100011: o_lut = 11'b01010100011;  // K.03.5, RDin = -1, RDout = -1
      10'b1010100100: o_lut = 11'b10101101011;  // K.04.5, RDin = -1, RDout = +1
      10'b1010100101: o_lut = 11'b01010100101;  // K.05.5, RDin = -1, RDout = -1
      10'b1010100110: o_lut = 11'b01010100110;  // K.06.5, RDin = -1, RDout = -1
      10'b1010100111: o_lut = 11'b01010000111;  // K.07.5, RDin = -1, RDout = -1
      10'b1010101000: o_lut = 11'b10101100111;  // K.08.5, RDin = -1, RDout = +1
      10'b1010101001: o_lut = 11'b01010101001;  // K.09.5, RDin = -1, RDout = -1
      10'b1010101010: o_lut = 11'b01010101010;  // K.10.5, RDin = -1, RDout = -1
      10'b1010101011: o_lut = 11'b01010001011;  // K.11.5, RDin = -1, RDout = -1
      10'b1010101100: o_lut = 11'b01010101100;  // K.12.5, RDin = -1, RDout = -1
      10'b1010101101: o_lut = 11'b01010001101;  // K.13.5, RDin = -1, RDout = -1
      10'b1010101110: o_lut = 11'b01010001110;  // K.14.5, RDin = -1, RDout = -1
      10'b1010101111: o_lut = 11'b10101111010;  // K.15.5, RDin = -1, RDout = +1
      10'b1010110000: o_lut = 11'b10101110110;  // K.16.5, RDin = -1, RDout = +1
      10'b1010110001: o_lut = 11'b01010110001;  // K.17.5, RDin = -1, RDout = -1
      10'b1010110010: o_lut = 11'b01010110010;  // K.18.5, RDin = -1, RDout = -1
      10'b1010110011: o_lut = 11'b01010010011;  // K.19.5, RDin = -1, RDout = -1
      10'b1010110100: o_lut = 11'b01010110100;  // K.20.5, RDin = -1, RDout = -1
      10'b1010110101: o_lut = 11'b01010010101;  // K.21.5, RDin = -1, RDout = -1
      10'b1010110110: o_lut = 11'b01010010110;  // K.22.5, RDin = -1, RDout = -1
      10'b1010110111: o_lut = 11'b10101010111;  // K.23.5, RDin = -1, RDout = +1
      10'b1010111000: o_lut = 11'b10101110011;  // K.24.5, RDin = -1, RDout = +1
      10'b1010111001: o_lut = 11'b01010011001;  // K.25.5, RDin = -1, RDout = -1
      10'b1010111010: o_lut = 11'b01010011010;  // K.26.5, RDin = -1, RDout = -1
      10'b1010111011: o_lut = 11'b10101011011;  // K.27.5, RDin = -1, RDout = +1
      10'b1010111100: o_lut = 11'b10101111100;  // K.28.5, RDin = -1, RDout = +1
      10'b1010111101: o_lut = 11'b10101011101;  // K.29.5, RDin = -1, RDout = +1
      10'b1010111110: o_lut = 11'b10101011110;  // K.30.5, RDin = -1, RDout = +1
      10'b1010111111: o_lut = 11'b10101110101;  // K.31.5, RDin = -1, RDout = +1
      10'b1011000000: o_lut = 11'b10110111001;  // K.00.6, RDin = -1, RDout = +1
      10'b1011000001: o_lut = 11'b10110101110;  // K.01.6, RDin = -1, RDout = +1
      10'b1011000010: o_lut = 11'b10110101101;  // K.02.6, RDin = -1, RDout = +1
      10'b1011000011: o_lut = 11'b01001100011;  // K.03.6, RDin = -1, RDout = -1
      10'b1011000100: o_lut = 11'b10110101011;  // K.04.6, RDin = -1, RDout = +1
      10'b1011000101: o_lut = 11'b01001100101;  // K.05.6, RDin = -1, RDout = -1
      10'b1011000110: o_lut = 11'b01001100110;  // K.06.6, RDin = -1, RDout = -1
      10'b1011000111: o_lut = 11'b01001000111;  // K.07.6, RDin = -1, RDout = -1
      10'b1011001000: o_lut = 11'b10110100111;  // K.08.6, RDin = -1, RDout = +1
      10'b1011001001: o_lut = 11'b01001101001;  // K.09.6, RDin = -1, RDout = -1
      10'b1011001010: o_lut = 11'b01001101010;  // K.10.6, RDin = -1, RDout = -1
      10'b1011001011: o_lut = 11'b01001001011;  // K.11.6, RDin = -1, RDout = -1
      10'b1011001100: o_lut = 11'b01001101100;  // K.12.6, RDin = -1, RDout = -1
      10'b1011001101: o_lut = 11'b01001001101;  // K.13.6, RDin = -1, RDout = -1
      10'b1011001110: o_lut = 11'b01001001110;  // K.14.6, RDin = -1, RDout = -1
      10'b1011001111: o_lut = 11'b10110111010;  // K.15.6, RDin = -1, RDout = +1
      10'b1011010000: o_lut = 11'b10110110110;  // K.16.6, RDin = -1, RDout = +1
      10'b1011010001: o_lut = 11'b01001110001;  // K.17.6, RDin = -1, RDout = -1
      10'b1011010010: o_lut = 11'b01001110010;  // K.18.6, RDin = -1, RDout = -1
      10'b1011010011: o_lut = 11'b01001010011;  // K.19.6, RDin = -1, RDout = -1
      10'b1011010100: o_lut = 11'b01001110100;  // K.20.6, RDin = -1, RDout = -1
      10'b1011010101: o_lut = 11'b01001010101;  // K.21.6, RDin = -1, RDout = -1
      10'b1011010110: o_lut = 11'b01001010110;  // K.22.6, RDin = -1, RDout = -1
      10'b1011010111: o_lut = 11'b10110010111;  // K.23.6, RDin = -1, RDout = +1
      10'b1011011000: o_lut = 11'b10110110011;  // K.24.6, RDin = -1, RDout = +1
      10'b1011011001: o_lut = 11'b01001011001;  // K.25.6, RDin = -1, RDout = -1
      10'b1011011010: o_lut = 11'b01001011010;  // K.26.6, RDin = -1, RDout = -1
      10'b1011011011: o_lut = 11'b10110011011;  // K.27.6, RDin = -1, RDout = +1
      10'b1011011100: o_lut = 11'b10110111100;  // K.28.6, RDin = -1, RDout = +1
      10'b1011011101: o_lut = 11'b10110011101;  // K.29.6, RDin = -1, RDout = +1
      10'b1011011110: o_lut = 11'b10110011110;  // K.30.6, RDin = -1, RDout = +1
      10'b1011011111: o_lut = 11'b10110110101;  // K.31.6, RDin = -1, RDout = +1
      10'b1011100000: o_lut = 11'b00001111001;  // K.00.7, RDin = -1, RDout = -1
      10'b1011100001: o_lut = 11'b00001101110;  // K.01.7, RDin = -1, RDout = -1
      10'b1011100010: o_lut = 11'b00001101101;  // K.02.7, RDin = -1, RDout = -1
      10'b1011100011: o_lut = 11'b11110100011;  // K.03.7, RDin = -1, RDout = +1
      10'b1011100100: o_lut = 11'b00001101011;  // K.04.7, RDin = -1, RDout = -1
      10'b1011100101: o_lut = 11'b11110100101;  // K.05.7, RDin = -1, RDout = +1
      10'b1011100110: o_lut = 11'b11110100110;  // K.06.7, RDin = -1, RDout = +1
      10'b1011100111: o_lut = 11'b11110000111;  // K.07.7, RDin = -1, RDout = +1
      10'b1011101000: o_lut = 11'b00001100111;  // K.08.7, RDin = -1, RDout = -1
      10'b1011101001: o_lut = 11'b11110101001;  // K.09.7, RDin = -1, RDout = +1
      10'b1011101010: o_lut = 11'b11110101010;  // K.10.7, RDin = -1, RDout = +1
      10'b1011101011: o_lut = 11'b11110001011;  // K.11.7, RDin = -1, RDout = +1
      10'b1011101100: o_lut = 11'b11110101100;  // K.12.7, RDin = -1, RDout = +1
      10'b1011101101: o_lut = 11'b11110001101;  // K.13.7, RDin = -1, RDout = +1
      10'b1011101110: o_lut = 11'b11110001110;  // K.14.7, RDin = -1, RDout = +1
      10'b1011101111: o_lut = 11'b00001111010;  // K.15.7, RDin = -1, RDout = -1
      10'b1011110000: o_lut = 11'b00001110110;  // K.16.7, RDin = -1, RDout = -1
      10'b1011110001: o_lut = 11'b11110110001;  // K.17.7, RDin = -1, RDout = +1
      10'b1011110010: o_lut = 11'b11110110010;  // K.18.7, RDin = -1, RDout = +1
      10'b1011110011: o_lut = 11'b11110010011;  // K.19.7, RDin = -1, RDout = +1
      10'b1011110100: o_lut = 11'b11110110100;  // K.20.7, RDin = -1, RDout = +1
      10'b1011110101: o_lut = 11'b11110010101;  // K.21.7, RDin = -1, RDout = +1
      10'b1011110110: o_lut = 11'b11110010110;  // K.22.7, RDin = -1, RDout = +1
      10'b1011110111: o_lut = 11'b00001010111;  // K.23.7, RDin = -1, RDout = -1
      10'b1011111000: o_lut = 11'b00001110011;  // K.24.7, RDin = -1, RDout = -1
      10'b1011111001: o_lut = 11'b11110011001;  // K.25.7, RDin = -1, RDout = +1
      10'b1011111010: o_lut = 11'b11110011010;  // K.26.7, RDin = -1, RDout = +1
      10'b1011111011: o_lut = 11'b00001011011;  // K.27.7, RDin = -1, RDout = -1
      10'b1011111100: o_lut = 11'b00001111100;  // K.28.7, RDin = -1, RDout = -1
      10'b1011111101: o_lut = 11'b00001011101;  // K.29.7, RDin = -1, RDout = -1
      10'b1011111110: o_lut = 11'b00001011110;  // K.30.7, RDin = -1, RDout = -1
      10'b1011111111: o_lut = 11'b00001110101;  // K.31.7, RDin = -1, RDout = -1
      10'b1100000000: o_lut = 11'b11101000110;  // K.00.0, RDin = +1, RDout = +1
      10'b1100000001: o_lut = 11'b11101010001;  // K.01.0, RDin = +1, RDout = +1
      10'b1100000010: o_lut = 11'b11101010010;  // K.02.0, RDin = +1, RDout = +1
      10'b1100000011: o_lut = 11'b00010100011;  // K.03.0, RDin = +1, RDout = -1
      10'b1100000100: o_lut = 11'b11101010100;  // K.04.0, RDin = +1, RDout = +1
      10'b1100000101: o_lut = 11'b00010100101;  // K.05.0, RDin = +1, RDout = -1
      10'b1100000110: o_lut = 11'b00010100110;  // K.06.0, RDin = +1, RDout = -1
      10'b1100000111: o_lut = 11'b00010111000;  // K.07.0, RDin = +1, RDout = -1
      10'b1100001000: o_lut = 11'b11101011000;  // K.08.0, RDin = +1, RDout = +1
      10'b1100001001: o_lut = 11'b00010101001;  // K.09.0, RDin = +1, RDout = -1
      10'b1100001010: o_lut = 11'b00010101010;  // K.10.0, RDin = +1, RDout = -1
      10'b1100001011: o_lut = 11'b00010001011;  // K.11.0, RDin = +1, RDout = -1
      10'b1100001100: o_lut = 11'b00010101100;  // K.12.0, RDin = +1, RDout = -1
      10'b1100001101: o_lut = 11'b00010001101;  // K.13.0, RDin = +1, RDout = -1
      10'b1100001110: o_lut = 11'b00010001110;  // K.14.0, RDin = +1, RDout = -1
      10'b1100001111: o_lut = 11'b11101000101;  // K.15.0, RDin = +1, RDout = +1
      10'b1100010000: o_lut = 11'b11101001001;  // K.16.0, RDin = +1, RDout = +1
      10'b1100010001: o_lut = 11'b00010110001;  // K.17.0, RDin = +1, RDout = -1
      10'b1100010010: o_lut = 11'b00010110010;  // K.18.0, RDin = +1, RDout = -1
      10'b1100010011: o_lut = 11'b00010010011;  // K.19.0, RDin = +1, RDout = -1
      10'b1100010100: o_lut = 11'b00010110100;  // K.20.0, RDin = +1, RDout = -1
      10'b1100010101: o_lut = 11'b00010010101;  // K.21.0, RDin = +1, RDout = -1
      10'b1100010110: o_lut = 11'b00010010110;  // K.22.0, RDin = +1, RDout = -1
      10'b1100010111: o_lut = 11'b11101101000;  // K.23.0, RDin = +1, RDout = +1
      10'b1100011000: o_lut = 11'b11101001100;  // K.24.0, RDin = +1, RDout = +1
      10'b1100011001: o_lut = 11'b00010011001;  // K.25.0, RDin = +1, RDout = -1
      10'b1100011010: o_lut = 11'b00010011010;  // K.26.0, RDin = +1, RDout = -1
      10'b1100011011: o_lut = 11'b11101100100;  // K.27.0, RDin = +1, RDout = +1
      10'b1100011100: o_lut = 11'b11101000011;  // K.28.0, RDin = +1, RDout = +1
      10'b1100011101: o_lut = 11'b11101100010;  // K.29.0, RDin = +1, RDout = +1
      10'b1100011110: o_lut = 11'b11101100001;  // K.30.0, RDin = +1, RDout = +1
      10'b1100011111: o_lut = 11'b11101001010;  // K.31.0, RDin = +1, RDout = +1
      10'b1100100000: o_lut = 11'b00110000110;  // K.00.1, RDin = +1, RDout = -1
      10'b1100100001: o_lut = 11'b00110010001;  // K.01.1, RDin = +1, RDout = -1
      10'b1100100010: o_lut = 11'b00110010010;  // K.02.1, RDin = +1, RDout = -1
      10'b1100100011: o_lut = 11'b11001100011;  // K.03.1, RDin = +1, RDout = +1
      10'b1100100100: o_lut = 11'b00110010100;  // K.04.1, RDin = +1, RDout = -1
      10'b1100100101: o_lut = 11'b11001100101;  // K.05.1, RDin = +1, RDout = +1
      10'b1100100110: o_lut = 11'b11001100110;  // K.06.1, RDin = +1, RDout = +1
      10'b1100100111: o_lut = 11'b11001111000;  // K.07.1, RDin = +1, RDout = +1
      10'b1100101000: o_lut = 11'b00110011000;  // K.08.1, RDin = +1, RDout = -1
      10'b1100101001: o_lut = 11'b11001101001;  // K.09.1, RDin = +1, RDout = +1
      10'b1100101010: o_lut = 11'b11001101010;  // K.10.1, RDin = +1, RDout = +1
      10'b1100101011: o_lut = 11'b11001001011;  // K.11.1, RDin = +1, RDout = +1
      10'b1100101100: o_lut = 11'b11001101100;  // K.12.1, RDin = +1, RDout = +1
      10'b1100101101: o_lut = 11'b11001001101;  // K.13.1, RDin = +1, RDout = +1
      10'b1100101110: o_lut = 11'b11001001110;  // K.14.1, RDin = +1, RDout = +1
      10'b1100101111: o_lut = 11'b00110000101;  // K.15.1, RDin = +1, RDout = -1
      10'b1100110000: o_lut = 11'b00110001001;  // K.16.1, RDin = +1, RDout = -1
      10'b1100110001: o_lut = 11'b11001110001;  // K.17.1, RDin = +1, RDout = +1
      10'b1100110010: o_lut = 11'b11001110010;  // K.18.1, RDin = +1, RDout = +1
      10'b1100110011: o_lut = 11'b11001010011;  // K.19.1, RDin = +1, RDout = +1
      10'b1100110100: o_lut = 11'b11001110100;  // K.20.1, RDin = +1, RDout = +1
      10'b1100110101: o_lut = 11'b11001010101;  // K.21.1, RDin = +1, RDout = +1
      10'b1100110110: o_lut = 11'b11001010110;  // K.22.1, RDin = +1, RDout = +1
      10'b1100110111: o_lut = 11'b00110101000;  // K.23.1, RDin = +1, RDout = -1
      10'b1100111000: o_lut = 11'b00110001100;  // K.24.1, RDin = +1, RDout = -1
      10'b1100111001: o_lut = 11'b11001011001;  // K.25.1, RDin = +1, RDout = +1
      10'b1100111010: o_lut = 11'b11001011010;  // K.26.1, RDin = +1, RDout = +1
      10'b1100111011: o_lut = 11'b00110100100;  // K.27.1, RDin = +1, RDout = -1
      10'b1100111100: o_lut = 11'b00110000011;  // K.28.1, RDin = +1, RDout = -1
      10'b1100111101: o_lut = 11'b00110100010;  // K.29.1, RDin = +1, RDout = -1
      10'b1100111110: o_lut = 11'b00110100001;  // K.30.1, RDin = +1, RDout = -1
      10'b1100111111: o_lut = 11'b00110001010;  // K.31.1, RDin = +1, RDout = -1
      10'b1101000000: o_lut = 11'b00101000110;  // K.00.2, RDin = +1, RDout = -1
      10'b1101000001: o_lut = 11'b00101010001;  // K.01.2, RDin = +1, RDout = -1
      10'b1101000010: o_lut = 11'b00101010010;  // K.02.2, RDin = +1, RDout = -1
      10'b1101000011: o_lut = 11'b11010100011;  // K.03.2, RDin = +1, RDout = +1
      10'b1101000100: o_lut = 11'b00101010100;  // K.04.2, RDin = +1, RDout = -1
      10'b1101000101: o_lut = 11'b11010100101;  // K.05.2, RDin = +1, RDout = +1
      10'b1101000110: o_lut = 11'b11010100110;  // K.06.2, RDin = +1, RDout = +1
      10'b1101000111: o_lut = 11'b11010111000;  // K.07.2, RDin = +1, RDout = +1
      10'b1101001000: o_lut = 11'b00101011000;  // K.08.2, RDin = +1, RDout = -1
      10'b1101001001: o_lut = 11'b11010101001;  // K.09.2, RDin = +1, RDout = +1
      10'b1101001010: o_lut = 11'b11010101010;  // K.10.2, RDin = +1, RDout = +1
      10'b1101001011: o_lut = 11'b11010001011;  // K.11.2, RDin = +1, RDout = +1
      10'b1101001100: o_lut = 11'b11010101100;  // K.12.2, RDin = +1, RDout = +1
      10'b1101001101: o_lut = 11'b11010001101;  // K.13.2, RDin = +1, RDout = +1
      10'b1101001110: o_lut = 11'b11010001110;  // K.14.2, RDin = +1, RDout = +1
      10'b1101001111: o_lut = 11'b00101000101;  // K.15.2, RDin = +1, RDout = -1
      10'b1101010000: o_lut = 11'b00101001001;  // K.16.2, RDin = +1, RDout = -1
      10'b1101010001: o_lut = 11'b11010110001;  // K.17.2, RDin = +1, RDout = +1
      10'b1101010010: o_lut = 11'b11010110010;  // K.18.2, RDin = +1, RDout = +1
      10'b1101010011: o_lut = 11'b11010010011;  // K.19.2, RDin = +1, RDout = +1
      10'b1101010100: o_lut = 11'b11010110100;  // K.20.2, RDin = +1, RDout = +1
      10'b1101010101: o_lut = 11'b11010010101;  // K.21.2, RDin = +1, RDout = +1
      10'b1101010110: o_lut = 11'b11010010110;  // K.22.2, RDin = +1, RDout = +1
      10'b1101010111: o_lut = 11'b00101101000;  // K.23.2, RDin = +1, RDout = -1
      10'b1101011000: o_lut = 11'b00101001100;  // K.24.2, RDin = +1, RDout = -1
      10'b1101011001: o_lut = 11'b11010011001;  // K.25.2, RDin = +1, RDout = +1
      10'b1101011010: o_lut = 11'b11010011010;  // K.26.2, RDin = +1, RDout = +1
      10'b1101011011: o_lut = 11'b00101100100;  // K.27.2, RDin = +1, RDout = -1
      10'b1101011100: o_lut = 11'b00101000011;  // K.28.2, RDin = +1, RDout = -1
      10'b1101011101: o_lut = 11'b00101100010;  // K.29.2, RDin = +1, RDout = -1
      10'b1101011110: o_lut = 11'b00101100001;  // K.30.2, RDin = +1, RDout = -1
      10'b1101011111: o_lut = 11'b00101001010;  // K.31.2, RDin = +1, RDout = -1
      10'b1101100000: o_lut = 11'b00011000110;  // K.00.3, RDin = +1, RDout = -1
      10'b1101100001: o_lut = 11'b00011010001;  // K.01.3, RDin = +1, RDout = -1
      10'b1101100010: o_lut = 11'b00011010010;  // K.02.3, RDin = +1, RDout = -1
      10'b1101100011: o_lut = 11'b11100100011;  // K.03.3, RDin = +1, RDout = +1
      10'b1101100100: o_lut = 11'b00011010100;  // K.04.3, RDin = +1, RDout = -1
      10'b1101100101: o_lut = 11'b11100100101;  // K.05.3, RDin = +1, RDout = +1
      10'b1101100110: o_lut = 11'b11100100110;  // K.06.3, RDin = +1, RDout = +1
      10'b1101100111: o_lut = 11'b11100111000;  // K.07.3, RDin = +1, RDout = +1
      10'b1101101000: o_lut = 11'b00011011000;  // K.08.3, RDin = +1, RDout = -1
      10'b1101101001: o_lut = 11'b11100101001;  // K.09.3, RDin = +1, RDout = +1
      10'b1101101010: o_lut = 11'b11100101010;  // K.10.3, RDin = +1, RDout = +1
      10'b1101101011: o_lut = 11'b11100001011;  // K.11.3, RDin = +1, RDout = +1
      10'b1101101100: o_lut = 11'b11100101100;  // K.12.3, RDin = +1, RDout = +1
      10'b1101101101: o_lut = 11'b11100001101;  // K.13.3, RDin = +1, RDout = +1
      10'b1101101110: o_lut = 11'b11100001110;  // K.14.3, RDin = +1, RDout = +1
      10'b1101101111: o_lut = 11'b00011000101;  // K.15.3, RDin = +1, RDout = -1
      10'b1101110000: o_lut = 11'b00011001001;  // K.16.3, RDin = +1, RDout = -1
      10'b1101110001: o_lut = 11'b11100110001;  // K.17.3, RDin = +1, RDout = +1
      10'b1101110010: o_lut = 11'b11100110010;  // K.18.3, RDin = +1, RDout = +1
      10'b1101110011: o_lut = 11'b11100010011;  // K.19.3, RDin = +1, RDout = +1
      10'b1101110100: o_lut = 11'b11100110100;  // K.20.3, RDin = +1, RDout = +1
      10'b1101110101: o_lut = 11'b11100010101;  // K.21.3, RDin = +1, RDout = +1
      10'b1101110110: o_lut = 11'b11100010110;  // K.22.3, RDin = +1, RDout = +1
      10'b1101110111: o_lut = 11'b00011101000;  // K.23.3, RDin = +1, RDout = -1
      10'b1101111000: o_lut = 11'b00011001100;  // K.24.3, RDin = +1, RDout = -1
      10'b1101111001: o_lut = 11'b11100011001;  // K.25.3, RDin = +1, RDout = +1
      10'b1101111010: o_lut = 11'b11100011010;  // K.26.3, RDin = +1, RDout = +1
      10'b1101111011: o_lut = 11'b00011100100;  // K.27.3, RDin = +1, RDout = -1
      10'b1101111100: o_lut = 11'b00011000011;  // K.28.3, RDin = +1, RDout = -1
      10'b1101111101: o_lut = 11'b00011100010;  // K.29.3, RDin = +1, RDout = -1
      10'b1101111110: o_lut = 11'b00011100001;  // K.30.3, RDin = +1, RDout = -1
      10'b1101111111: o_lut = 11'b00011001010;  // K.31.3, RDin = +1, RDout = -1
      10'b1110000000: o_lut = 11'b11011000110;  // K.00.4, RDin = +1, RDout = +1
      10'b1110000001: o_lut = 11'b11011010001;  // K.01.4, RDin = +1, RDout = +1
      10'b1110000010: o_lut = 11'b11011010010;  // K.02.4, RDin = +1, RDout = +1
      10'b1110000011: o_lut = 11'b00100100011;  // K.03.4, RDin = +1, RDout = -1
      10'b1110000100: o_lut = 11'b11011010100;  // K.04.4, RDin = +1, RDout = +1
      10'b1110000101: o_lut = 11'b00100100101;  // K.05.4, RDin = +1, RDout = -1
      10'b1110000110: o_lut = 11'b00100100110;  // K.06.4, RDin = +1, RDout = -1
      10'b1110000111: o_lut = 11'b00100111000;  // K.07.4, RDin = +1, RDout = -1
      10'b1110001000: o_lut = 11'b11011011000;  // K.08.4, RDin = +1, RDout = +1
      10'b1110001001: o_lut = 11'b00100101001;  // K.09.4, RDin = +1, RDout = -1
      10'b1110001010: o_lut = 11'b00100101010;  // K.10.4, RDin = +1, RDout = -1
      10'b1110001011: o_lut = 11'b00100001011;  // K.11.4, RDin = +1, RDout = -1
      10'b1110001100: o_lut = 11'b00100101100;  // K.12.4, RDin = +1, RDout = -1
      10'b1110001101: o_lut = 11'b00100001101;  // K.13.4, RDin = +1, RDout = -1
      10'b1110001110: o_lut = 11'b00100001110;  // K.14.4, RDin = +1, RDout = -1
      10'b1110001111: o_lut = 11'b11011000101;  // K.15.4, RDin = +1, RDout = +1
      10'b1110010000: o_lut = 11'b11011001001;  // K.16.4, RDin = +1, RDout = +1
      10'b1110010001: o_lut = 11'b00100110001;  // K.17.4, RDin = +1, RDout = -1
      10'b1110010010: o_lut = 11'b00100110010;  // K.18.4, RDin = +1, RDout = -1
      10'b1110010011: o_lut = 11'b00100010011;  // K.19.4, RDin = +1, RDout = -1
      10'b1110010100: o_lut = 11'b00100110100;  // K.20.4, RDin = +1, RDout = -1
      10'b1110010101: o_lut = 11'b00100010101;  // K.21.4, RDin = +1, RDout = -1
      10'b1110010110: o_lut = 11'b00100010110;  // K.22.4, RDin = +1, RDout = -1
      10'b1110010111: o_lut = 11'b11011101000;  // K.23.4, RDin = +1, RDout = +1
      10'b1110011000: o_lut = 11'b11011001100;  // K.24.4, RDin = +1, RDout = +1
      10'b1110011001: o_lut = 11'b00100011001;  // K.25.4, RDin = +1, RDout = -1
      10'b1110011010: o_lut = 11'b00100011010;  // K.26.4, RDin = +1, RDout = -1
      10'b1110011011: o_lut = 11'b11011100100;  // K.27.4, RDin = +1, RDout = +1
      10'b1110011100: o_lut = 11'b11011000011;  // K.28.4, RDin = +1, RDout = +1
      10'b1110011101: o_lut = 11'b11011100010;  // K.29.4, RDin = +1, RDout = +1
      10'b1110011110: o_lut = 11'b11011100001;  // K.30.4, RDin = +1, RDout = +1
      10'b1110011111: o_lut = 11'b11011001010;  // K.31.4, RDin = +1, RDout = +1
      10'b1110100000: o_lut = 11'b01010000110;  // K.00.5, RDin = +1, RDout = -1
      10'b1110100001: o_lut = 11'b01010010001;  // K.01.5, RDin = +1, RDout = -1
      10'b1110100010: o_lut = 11'b01010010010;  // K.02.5, RDin = +1, RDout = -1
      10'b1110100011: o_lut = 11'b10101100011;  // K.03.5, RDin = +1, RDout = +1
      10'b1110100100: o_lut = 11'b01010010100;  // K.04.5, RDin = +1, RDout = -1
      10'b1110100101: o_lut = 11'b10101100101;  // K.05.5, RDin = +1, RDout = +1
      10'b1110100110: o_lut = 11'b10101100110;  // K.06.5, RDin = +1, RDout = +1
      10'b1110100111: o_lut = 11'b10101111000;  // K.07.5, RDin = +1, RDout = +1
      10'b1110101000: o_lut = 11'b01010011000;  // K.08.5, RDin = +1, RDout = -1
      10'b1110101001: o_lut = 11'b10101101001;  // K.09.5, RDin = +1, RDout = +1
      10'b1110101010: o_lut = 11'b10101101010;  // K.10.5, RDin = +1, RDout = +1
      10'b1110101011: o_lut = 11'b10101001011;  // K.11.5, RDin = +1, RDout = +1
      10'b1110101100: o_lut = 11'b10101101100;  // K.12.5, RDin = +1, RDout = +1
      10'b1110101101: o_lut = 11'b10101001101;  // K.13.5, RDin = +1, RDout = +1
      10'b1110101110: o_lut = 11'b10101001110;  // K.14.5, RDin = +1, RDout = +1
      10'b1110101111: o_lut = 11'b01010000101;  // K.15.5, RDin = +1, RDout = -1
      10'b1110110000: o_lut = 11'b01010001001;  // K.16.5, RDin = +1, RDout = -1
      10'b1110110001: o_lut = 11'b10101110001;  // K.17.5, RDin = +1, RDout = +1
      10'b1110110010: o_lut = 11'b10101110010;  // K.18.5, RDin = +1, RDout = +1
      10'b1110110011: o_lut = 11'b10101010011;  // K.19.5, RDin = +1, RDout = +1
      10'b1110110100: o_lut = 11'b10101110100;  // K.20.5, RDin = +1, RDout = +1
      10'b1110110101: o_lut = 11'b10101010101;  // K.21.5, RDin = +1, RDout = +1
      10'b1110110110: o_lut = 11'b10101010110;  // K.22.5, RDin = +1, RDout = +1
      10'b1110110111: o_lut = 11'b01010101000;  // K.23.5, RDin = +1, RDout = -1
      10'b1110111000: o_lut = 11'b01010001100;  // K.24.5, RDin = +1, RDout = -1
      10'b1110111001: o_lut = 11'b10101011001;  // K.25.5, RDin = +1, RDout = +1
      10'b1110111010: o_lut = 11'b10101011010;  // K.26.5, RDin = +1, RDout = +1
      10'b1110111011: o_lut = 11'b01010100100;  // K.27.5, RDin = +1, RDout = -1
      10'b1110111100: o_lut = 11'b01010000011;  // K.28.5, RDin = +1, RDout = -1
      10'b1110111101: o_lut = 11'b01010100010;  // K.29.5, RDin = +1, RDout = -1
      10'b1110111110: o_lut = 11'b01010100001;  // K.30.5, RDin = +1, RDout = -1
      10'b1110111111: o_lut = 11'b01010001010;  // K.31.5, RDin = +1, RDout = -1
      10'b1111000000: o_lut = 11'b01001000110;  // K.00.6, RDin = +1, RDout = -1
      10'b1111000001: o_lut = 11'b01001010001;  // K.01.6, RDin = +1, RDout = -1
      10'b1111000010: o_lut = 11'b01001010010;  // K.02.6, RDin = +1, RDout = -1
      10'b1111000011: o_lut = 11'b10110100011;  // K.03.6, RDin = +1, RDout = +1
      10'b1111000100: o_lut = 11'b01001010100;  // K.04.6, RDin = +1, RDout = -1
      10'b1111000101: o_lut = 11'b10110100101;  // K.05.6, RDin = +1, RDout = +1
      10'b1111000110: o_lut = 11'b10110100110;  // K.06.6, RDin = +1, RDout = +1
      10'b1111000111: o_lut = 11'b10110111000;  // K.07.6, RDin = +1, RDout = +1
      10'b1111001000: o_lut = 11'b01001011000;  // K.08.6, RDin = +1, RDout = -1
      10'b1111001001: o_lut = 11'b10110101001;  // K.09.6, RDin = +1, RDout = +1
      10'b1111001010: o_lut = 11'b10110101010;  // K.10.6, RDin = +1, RDout = +1
      10'b1111001011: o_lut = 11'b10110001011;  // K.11.6, RDin = +1, RDout = +1
      10'b1111001100: o_lut = 11'b10110101100;  // K.12.6, RDin = +1, RDout = +1
      10'b1111001101: o_lut = 11'b10110001101;  // K.13.6, RDin = +1, RDout = +1
      10'b1111001110: o_lut = 11'b10110001110;  // K.14.6, RDin = +1, RDout = +1
      10'b1111001111: o_lut = 11'b01001000101;  // K.15.6, RDin = +1, RDout = -1
      10'b1111010000: o_lut = 11'b01001001001;  // K.16.6, RDin = +1, RDout = -1
      10'b1111010001: o_lut = 11'b10110110001;  // K.17.6, RDin = +1, RDout = +1
      10'b1111010010: o_lut = 11'b10110110010;  // K.18.6, RDin = +1, RDout = +1
      10'b1111010011: o_lut = 11'b10110010011;  // K.19.6, RDin = +1, RDout = +1
      10'b1111010100: o_lut = 11'b10110110100;  // K.20.6, RDin = +1, RDout = +1
      10'b1111010101: o_lut = 11'b10110010101;  // K.21.6, RDin = +1, RDout = +1
      10'b1111010110: o_lut = 11'b10110010110;  // K.22.6, RDin = +1, RDout = +1
      10'b1111010111: o_lut = 11'b01001101000;  // K.23.6, RDin = +1, RDout = -1
      10'b1111011000: o_lut = 11'b01001001100;  // K.24.6, RDin = +1, RDout = -1
      10'b1111011001: o_lut = 11'b10110011001;  // K.25.6, RDin = +1, RDout = +1
      10'b1111011010: o_lut = 11'b10110011010;  // K.26.6, RDin = +1, RDout = +1
      10'b1111011011: o_lut = 11'b01001100100;  // K.27.6, RDin = +1, RDout = -1
      10'b1111011100: o_lut = 11'b01001000011;  // K.28.6, RDin = +1, RDout = -1
      10'b1111011101: o_lut = 11'b01001100010;  // K.29.6, RDin = +1, RDout = -1
      10'b1111011110: o_lut = 11'b01001100001;  // K.30.6, RDin = +1, RDout = -1
      10'b1111011111: o_lut = 11'b01001001010;  // K.31.6, RDin = +1, RDout = -1
      10'b1111100000: o_lut = 11'b11110000110;  // K.00.7, RDin = +1, RDout = +1
      10'b1111100001: o_lut = 11'b11110010001;  // K.01.7, RDin = +1, RDout = +1
      10'b1111100010: o_lut = 11'b11110010010;  // K.02.7, RDin = +1, RDout = +1
      10'b1111100011: o_lut = 11'b00001100011;  // K.03.7, RDin = +1, RDout = -1
      10'b1111100100: o_lut = 11'b11110010100;  // K.04.7, RDin = +1, RDout = +1
      10'b1111100101: o_lut = 11'b00001100101;  // K.05.7, RDin = +1, RDout = -1
      10'b1111100110: o_lut = 11'b00001100110;  // K.06.7, RDin = +1, RDout = -1
      10'b1111100111: o_lut = 11'b00001111000;  // K.07.7, RDin = +1, RDout = -1
      10'b1111101000: o_lut = 11'b11110011000;  // K.08.7, RDin = +1, RDout = +1
      10'b1111101001: o_lut = 11'b00001101001;  // K.09.7, RDin = +1, RDout = -1
      10'b1111101010: o_lut = 11'b00001101010;  // K.10.7, RDin = +1, RDout = -1
      10'b1111101011: o_lut = 11'b00001001011;  // K.11.7, RDin = +1, RDout = -1
      10'b1111101100: o_lut = 11'b00001101100;  // K.12.7, RDin = +1, RDout = -1
      10'b1111101101: o_lut = 11'b00001001101;  // K.13.7, RDin = +1, RDout = -1
      10'b1111101110: o_lut = 11'b00001001110;  // K.14.7, RDin = +1, RDout = -1
      10'b1111101111: o_lut = 11'b11110000101;  // K.15.7, RDin = +1, RDout = +1
      10'b1111110000: o_lut = 11'b11110001001;  // K.16.7, RDin = +1, RDout = +1
      10'b1111110001: o_lut = 11'b00001110001;  // K.17.7, RDin = +1, RDout = -1
      10'b1111110010: o_lut = 11'b00001110010;  // K.18.7, RDin = +1, RDout = -1
      10'b1111110011: o_lut = 11'b00001010011;  // K.19.7, RDin = +1, RDout = -1
      10'b1111110100: o_lut = 11'b00001110100;  // K.20.7, RDin = +1, RDout = -1
      10'b1111110101: o_lut = 11'b00001010101;  // K.21.7, RDin = +1, RDout = -1
      10'b1111110110: o_lut = 11'b00001010110;  // K.22.7, RDin = +1, RDout = -1
      10'b1111110111: o_lut = 11'b11110101000;  // K.23.7, RDin = +1, RDout = +1
      10'b1111111000: o_lut = 11'b11110001100;  // K.24.7, RDin = +1, RDout = +1
      10'b1111111001: o_lut = 11'b00001011001;  // K.25.7, RDin = +1, RDout = -1
      10'b1111111010: o_lut = 11'b00001011010;  // K.26.7, RDin = +1, RDout = -1
      10'b1111111011: o_lut = 11'b11110100100;  // K.27.7, RDin = +1, RDout = +1
      10'b1111111100: o_lut = 11'b11110000011;  // K.28.7, RDin = +1, RDout = +1
      10'b1111111101: o_lut = 11'b11110100010;  // K.29.7, RDin = +1, RDout = +1
      10'b1111111110: o_lut = 11'b11110100001;  // K.30.7, RDin = +1, RDout = +1
      10'b1111111111: o_lut = 11'b11110001010;  // K.31.7, RDin = +1, RDout = +1
      default:        o_lut = 11'b11110001010;  // K.31.7, RDin = +1, RDout = +1
    endcase
  end

endmodule
